-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM80 is
	port(
		CE_n	: in std_logic;
		OE_n	: in std_logic;
		A	: in std_logic_vector(14 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end ROM80;

architecture rtl of ROM80 is
	subtype ROM_WORD is std_logic_vector(7 downto 0);
	type ROM_TABLE is array(0 to 8191) of ROM_WORD;
	constant ROM: ROM_TABLE := ROM_TABLE'(
		"11110011",	-- 0x0000
		"00011000",	-- 0x0001
		"00111010",	-- 0x0002
		"00000000",	-- 0x0003
		"00000000",	-- 0x0004
		"00000000",	-- 0x0005
		"00000000",	-- 0x0006
		"00000000",	-- 0x0007
		"11000101",	-- 0x0008
		"11100101",	-- 0x0009
		"11011101",	-- 0x000A
		"11100101",	-- 0x000B
		"11100001",	-- 0x000C
		"00101001",	-- 0x000D
		"00000001",	-- 0x000E
		"00011101",	-- 0x000F
		"00000000",	-- 0x0010
		"00001001",	-- 0x0011
		"01001110",	-- 0x0012
		"00100011",	-- 0x0013
		"01000110",	-- 0x0014
		"00101011",	-- 0x0015
		"11000101",	-- 0x0016
		"11011101",	-- 0x0017
		"11100001",	-- 0x0018
		"11100001",	-- 0x0019
		"11000001",	-- 0x001A
		"11011101",	-- 0x001B
		"11101001",	-- 0x001C
		"00110101",	-- 0x001D
		"00001101",	-- 0x001E
		"10010001",	-- 0x001F
		"00001010",	-- 0x0020
		"10100101",	-- 0x0021
		"00001010",	-- 0x0022
		"10111001",	-- 0x0023
		"00001010",	-- 0x0024
		"11010100",	-- 0x0025
		"00001010",	-- 0x0026
		"11100001",	-- 0x0027
		"00001010",	-- 0x0028
		"01100011",	-- 0x0029
		"00001011",	-- 0x002A
		"01101001",	-- 0x002B
		"00001011",	-- 0x002C
		"11000010",	-- 0x002D
		"00001010",	-- 0x002E
		"00010111",	-- 0x002F
		"00001011",	-- 0x0030
		"01111010",	-- 0x0031
		"00001101",	-- 0x0032
		"10100101",	-- 0x0033
		"00001110",	-- 0x0034
		"00110101",	-- 0x0035
		"00010000",	-- 0x0036
		"10000110",	-- 0x0037
		"00010001",	-- 0x0038
		"01100001",	-- 0x0039
		"00010011",	-- 0x003A
		"01011001",	-- 0x003B
		"00010110",	-- 0x003C
		"00110001",	-- 0x003D
		"01001011",	-- 0x003E
		"11111011",	-- 0x003F
		"00111110",	-- 0x0040
		"10000000",	-- 0x0041
		"11010011",	-- 0x0042
		"00000011",	-- 0x0043
		"00111110",	-- 0x0044
		"00001100",	-- 0x0045
		"11010011",	-- 0x0046
		"00000000",	-- 0x0047
		"10101111",	-- 0x0048
		"11010011",	-- 0x0049
		"00000001",	-- 0x004A
		"00111110",	-- 0x004B
		"00000011",	-- 0x004C
		"11010011",	-- 0x004D
		"00000011",	-- 0x004E
		"00100001",	-- 0x004F
		"01010011",	-- 0x0050
		"00000001",	-- 0x0051
		"11001101",	-- 0x0052
		"01101001",	-- 0x0053
		"00001011",	-- 0x0054
		"00111010",	-- 0x0055
		"01001100",	-- 0x0056
		"11111011",	-- 0x0057
		"11111110",	-- 0x0058
		"10101010",	-- 0x0059
		"00101000",	-- 0x005A
		"00011000",	-- 0x005B
		"00100001",	-- 0x005C
		"00000100",	-- 0x005D
		"00000010",	-- 0x005E
		"11001101",	-- 0x005F
		"01101001",	-- 0x0060
		"00001011",	-- 0x0061
		"00100001",	-- 0x0062
		"00000000",	-- 0x0063
		"10000000",	-- 0x0064
		"01010100",	-- 0x0065
		"01011101",	-- 0x0066
		"00010011",	-- 0x0067
		"00000001",	-- 0x0068
		"11111111",	-- 0x0069
		"01111111",	-- 0x006A
		"00110110",	-- 0x006B
		"00000000",	-- 0x006C
		"11101101",	-- 0x006D
		"10110000",	-- 0x006E
		"00100001",	-- 0x006F
		"01001100",	-- 0x0070
		"11111011",	-- 0x0071
		"00110110",	-- 0x0072
		"10101010",	-- 0x0073
		"00100001",	-- 0x0074
		"10010111",	-- 0x0075
		"00000001",	-- 0x0076
		"11001101",	-- 0x0077
		"01101001",	-- 0x0078
		"00001011",	-- 0x0079
		"11001101",	-- 0x007A
		"00100011",	-- 0x007B
		"00000010",	-- 0x007C
		"11111110",	-- 0x007D
		"01000011",	-- 0x007E
		"00100000",	-- 0x007F
		"00100010",	-- 0x0080
		"00100001",	-- 0x0081
		"10011101",	-- 0x0082
		"00000001",	-- 0x0083
		"11001101",	-- 0x0084
		"01101001",	-- 0x0085
		"00001011",	-- 0x0086
		"11001101",	-- 0x0087
		"00100011",	-- 0x0088
		"00000010",	-- 0x0089
		"11111110",	-- 0x008A
		"01000011",	-- 0x008B
		"11001010",	-- 0x008C
		"00110101",	-- 0x008D
		"00001101",	-- 0x008E
		"11111110",	-- 0x008F
		"01010111",	-- 0x0090
		"11001010",	-- 0x0091
		"00111010",	-- 0x0092
		"00001101",	-- 0x0093
		"11111110",	-- 0x0094
		"01010011",	-- 0x0095
		"11001010",	-- 0x0096
		"01100001",	-- 0x0097
		"00001010",	-- 0x0098
		"11111110",	-- 0x0099
		"01001001",	-- 0x009A
		"11001100",	-- 0x009B
		"10110101",	-- 0x009C
		"00000111",	-- 0x009D
		"00101000",	-- 0x009E
		"11010100",	-- 0x009F
		"11000011",	-- 0x00A0
		"01000111",	-- 0x00A1
		"00000001",	-- 0x00A2
		"11111110",	-- 0x00A3
		"01000100",	-- 0x00A4
		"00100000",	-- 0x00A5
		"00100111",	-- 0x00A6
		"00100001",	-- 0x00A7
		"10100110",	-- 0x00A8
		"00000001",	-- 0x00A9
		"11001101",	-- 0x00AA
		"01101001",	-- 0x00AB
		"00001011",	-- 0x00AC
		"11001101",	-- 0x00AD
		"00100011",	-- 0x00AE
		"00000010",	-- 0x00AF
		"11111110",	-- 0x00B0
		"01001001",	-- 0x00B1
		"11001100",	-- 0x00B2
		"10001000",	-- 0x00B3
		"00000010",	-- 0x00B4
		"00101000",	-- 0x00B5
		"10111101",	-- 0x00B6
		"11111110",	-- 0x00B7
		"01001101",	-- 0x00B8
		"11001100",	-- 0x00B9
		"00010111",	-- 0x00BA
		"00001001",	-- 0x00BB
		"00101000",	-- 0x00BC
		"10110110",	-- 0x00BD
		"11111110",	-- 0x00BE
		"01010100",	-- 0x00BF
		"11001100",	-- 0x00C0
		"10110100",	-- 0x00C1
		"00000010",	-- 0x00C2
		"00101000",	-- 0x00C3
		"10101111",	-- 0x00C4
		"11111110",	-- 0x00C5
		"01010101",	-- 0x00C6
		"11001100",	-- 0x00C7
		"01111011",	-- 0x00C8
		"00001010",	-- 0x00C9
		"00101000",	-- 0x00CA
		"10101000",	-- 0x00CB
		"00011000",	-- 0x00CC
		"01111001",	-- 0x00CD
		"11111110",	-- 0x00CE
		"01000110",	-- 0x00CF
		"00100000",	-- 0x00D0
		"00100000",	-- 0x00D1
		"00100001",	-- 0x00D2
		"10101100",	-- 0x00D3
		"00000001",	-- 0x00D4
		"11001101",	-- 0x00D5
		"01101001",	-- 0x00D6
		"00001011",	-- 0x00D7
		"11001101",	-- 0x00D8
		"00100011",	-- 0x00D9
		"00000010",	-- 0x00DA
		"11111110",	-- 0x00DB
		"01000011",	-- 0x00DC
		"11001100",	-- 0x00DD
		"00110100",	-- 0x00DE
		"00000010",	-- 0x00DF
		"00101000",	-- 0x00E0
		"10010010",	-- 0x00E1
		"11111110",	-- 0x00E2
		"01000100",	-- 0x00E3
		"11001100",	-- 0x00E4
		"01110000",	-- 0x00E5
		"00000010",	-- 0x00E6
		"00101000",	-- 0x00E7
		"10001011",	-- 0x00E8
		"11111110",	-- 0x00E9
		"01001100",	-- 0x00EA
		"11001100",	-- 0x00EB
		"01111001",	-- 0x00EC
		"00001000",	-- 0x00ED
		"00101000",	-- 0x00EE
		"10000100",	-- 0x00EF
		"00011000",	-- 0x00F0
		"01010101",	-- 0x00F1
		"11111110",	-- 0x00F2
		"01001000",	-- 0x00F3
		"11001100",	-- 0x00F4
		"00110001",	-- 0x00F5
		"00000101",	-- 0x00F6
		"11001010",	-- 0x00F7
		"01110100",	-- 0x00F8
		"00000000",	-- 0x00F9
		"11111110",	-- 0x00FA
		"01001101",	-- 0x00FB
		"11000010",	-- 0x00FC
		"01000010",	-- 0x00FD
		"00000001",	-- 0x00FE
		"00100001",	-- 0x00FF
		"10110010",	-- 0x0100
		"00000001",	-- 0x0101
		"11001101",	-- 0x0102
		"01101001",	-- 0x0103
		"00001011",	-- 0x0104
		"11001101",	-- 0x0105
		"00100011",	-- 0x0106
		"00000010",	-- 0x0107
		"11111110",	-- 0x0108
		"01000100",	-- 0x0109
		"11001100",	-- 0x010A
		"11000001",	-- 0x010B
		"00000011",	-- 0x010C
		"11001010",	-- 0x010D
		"01110100",	-- 0x010E
		"00000000",	-- 0x010F
		"11111110",	-- 0x0110
		"01000101",	-- 0x0111
		"11001100",	-- 0x0112
		"00110111",	-- 0x0113
		"00000100",	-- 0x0114
		"11001010",	-- 0x0115
		"01110100",	-- 0x0116
		"00000000",	-- 0x0117
		"11111110",	-- 0x0118
		"01000110",	-- 0x0119
		"11001100",	-- 0x011A
		"10001010",	-- 0x011B
		"00000100",	-- 0x011C
		"11001010",	-- 0x011D
		"01110100",	-- 0x011E
		"00000000",	-- 0x011F
		"11111110",	-- 0x0120
		"01001001",	-- 0x0121
		"11001100",	-- 0x0122
		"00000001",	-- 0x0123
		"00000111",	-- 0x0124
		"11001010",	-- 0x0125
		"01110100",	-- 0x0126
		"00000000",	-- 0x0127
		"11111110",	-- 0x0128
		"01001100",	-- 0x0129
		"11001100",	-- 0x012A
		"11001011",	-- 0x012B
		"00000111",	-- 0x012C
		"11001010",	-- 0x012D
		"01110100",	-- 0x012E
		"00000000",	-- 0x012F
		"11111110",	-- 0x0130
		"01001101",	-- 0x0131
		"11001100",	-- 0x0132
		"00101101",	-- 0x0133
		"00001001",	-- 0x0134
		"11001010",	-- 0x0135
		"01110100",	-- 0x0136
		"00000000",	-- 0x0137
		"11111110",	-- 0x0138
		"01010010",	-- 0x0139
		"11001100",	-- 0x013A
		"10100101",	-- 0x013B
		"00001001",	-- 0x013C
		"11001010",	-- 0x013D
		"01110100",	-- 0x013E
		"00000000",	-- 0x013F
		"00011000",	-- 0x0140
		"00000101",	-- 0x0141
		"00100001",	-- 0x0142
		"11100000",	-- 0x0143
		"00000001",	-- 0x0144
		"00011000",	-- 0x0145
		"00000011",	-- 0x0146
		"00100001",	-- 0x0147
		"10111010",	-- 0x0148
		"00000001",	-- 0x0149
		"11001101",	-- 0x014A
		"01100011",	-- 0x014B
		"00001011",	-- 0x014C
		"11001101",	-- 0x014D
		"01101001",	-- 0x014E
		"00001011",	-- 0x014F
		"11000011",	-- 0x0150
		"01110100",	-- 0x0151
		"00000000",	-- 0x0152
		"00001101",	-- 0x0153
		"00001010",	-- 0x0154
		"00001101",	-- 0x0155
		"00001010",	-- 0x0156
		"01010011",	-- 0x0157
		"01101001",	-- 0x0158
		"01101101",	-- 0x0159
		"01110000",	-- 0x015A
		"01101100",	-- 0x015B
		"01100101",	-- 0x015C
		"00100000",	-- 0x015D
		"01011010",	-- 0x015E
		"00111000",	-- 0x015F
		"00110000",	-- 0x0160
		"00101101",	-- 0x0161
		"01101101",	-- 0x0162
		"01101111",	-- 0x0163
		"01101110",	-- 0x0164
		"01101001",	-- 0x0165
		"01110100",	-- 0x0166
		"01101111",	-- 0x0167
		"01110010",	-- 0x0168
		"00100000",	-- 0x0169
		"00101101",	-- 0x016A
		"00100000",	-- 0x016B
		"01010110",	-- 0x016C
		"00100000",	-- 0x016D
		"00110000",	-- 0x016E
		"00101110",	-- 0x016F
		"00111000",	-- 0x0170
		"00100000",	-- 0x0171
		"00101000",	-- 0x0172
		"01000010",	-- 0x0173
		"00101110",	-- 0x0174
		"00100000",	-- 0x0175
		"01010101",	-- 0x0176
		"01101100",	-- 0x0177
		"01101101",	-- 0x0178
		"01100001",	-- 0x0179
		"01101110",	-- 0x017A
		"01101110",	-- 0x017B
		"00101100",	-- 0x017C
		"00100000",	-- 0x017D
		"01010011",	-- 0x017E
		"01100101",	-- 0x017F
		"01110000",	-- 0x0180
		"00101110",	-- 0x0181
		"00100000",	-- 0x0182
		"00110010",	-- 0x0183
		"00110000",	-- 0x0184
		"00110001",	-- 0x0185
		"00110001",	-- 0x0186
		"00100000",	-- 0x0187
		"00101101",	-- 0x0188
		"00100000",	-- 0x0189
		"01001010",	-- 0x018A
		"01100001",	-- 0x018B
		"01101110",	-- 0x018C
		"00101110",	-- 0x018D
		"00100000",	-- 0x018E
		"00110010",	-- 0x018F
		"00110000",	-- 0x0190
		"00110001",	-- 0x0191
		"00110010",	-- 0x0192
		"00101001",	-- 0x0193
		"00001101",	-- 0x0194
		"00001010",	-- 0x0195
		"00000000",	-- 0x0196
		"00001101",	-- 0x0197
		"00001010",	-- 0x0198
		"01011010",	-- 0x0199
		"00111110",	-- 0x019A
		"00100000",	-- 0x019B
		"00000000",	-- 0x019C
		"01000011",	-- 0x019D
		"01001111",	-- 0x019E
		"01001110",	-- 0x019F
		"01010100",	-- 0x01A0
		"01010010",	-- 0x01A1
		"01001111",	-- 0x01A2
		"01001100",	-- 0x01A3
		"00101111",	-- 0x01A4
		"00000000",	-- 0x01A5
		"01000100",	-- 0x01A6
		"01001001",	-- 0x01A7
		"01010011",	-- 0x01A8
		"01001011",	-- 0x01A9
		"00101111",	-- 0x01AA
		"00000000",	-- 0x01AB
		"01000110",	-- 0x01AC
		"01001001",	-- 0x01AD
		"01001100",	-- 0x01AE
		"01000101",	-- 0x01AF
		"00101111",	-- 0x01B0
		"00000000",	-- 0x01B1
		"01001101",	-- 0x01B2
		"01000101",	-- 0x01B3
		"01001101",	-- 0x01B4
		"01001111",	-- 0x01B5
		"01010010",	-- 0x01B6
		"01011001",	-- 0x01B7
		"00101111",	-- 0x01B8
		"00000000",	-- 0x01B9
		"00111010",	-- 0x01BA
		"00100000",	-- 0x01BB
		"01010011",	-- 0x01BC
		"01111001",	-- 0x01BD
		"01101110",	-- 0x01BE
		"01110100",	-- 0x01BF
		"01100001",	-- 0x01C0
		"01111000",	-- 0x01C1
		"00100000",	-- 0x01C2
		"01100101",	-- 0x01C3
		"01110010",	-- 0x01C4
		"01110010",	-- 0x01C5
		"01101111",	-- 0x01C6
		"01110010",	-- 0x01C7
		"00100000",	-- 0x01C8
		"00101101",	-- 0x01C9
		"00100000",	-- 0x01CA
		"01100011",	-- 0x01CB
		"01101111",	-- 0x01CC
		"01101101",	-- 0x01CD
		"01101101",	-- 0x01CE
		"01100001",	-- 0x01CF
		"01101110",	-- 0x01D0
		"01100100",	-- 0x01D1
		"00100000",	-- 0x01D2
		"01101110",	-- 0x01D3
		"01101111",	-- 0x01D4
		"01110100",	-- 0x01D5
		"00100000",	-- 0x01D6
		"01100110",	-- 0x01D7
		"01101111",	-- 0x01D8
		"01110101",	-- 0x01D9
		"01101110",	-- 0x01DA
		"01100100",	-- 0x01DB
		"00100001",	-- 0x01DC
		"00001101",	-- 0x01DD
		"00001010",	-- 0x01DE
		"00000000",	-- 0x01DF
		"00111010",	-- 0x01E0
		"00100000",	-- 0x01E1
		"01010011",	-- 0x01E2
		"01111001",	-- 0x01E3
		"01101110",	-- 0x01E4
		"01110100",	-- 0x01E5
		"01100001",	-- 0x01E6
		"01111000",	-- 0x01E7
		"00100000",	-- 0x01E8
		"01100101",	-- 0x01E9
		"01110010",	-- 0x01EA
		"01110010",	-- 0x01EB
		"01101111",	-- 0x01EC
		"01110010",	-- 0x01ED
		"00100000",	-- 0x01EE
		"00101101",	-- 0x01EF
		"00100000",	-- 0x01F0
		"01100111",	-- 0x01F1
		"01110010",	-- 0x01F2
		"01101111",	-- 0x01F3
		"01110101",	-- 0x01F4
		"01110000",	-- 0x01F5
		"00100000",	-- 0x01F6
		"01101110",	-- 0x01F7
		"01101111",	-- 0x01F8
		"01110100",	-- 0x01F9
		"00100000",	-- 0x01FA
		"01100110",	-- 0x01FB
		"01101111",	-- 0x01FC
		"01110101",	-- 0x01FD
		"01101110",	-- 0x01FE
		"01100100",	-- 0x01FF
		"00100001",	-- 0x0200
		"00001101",	-- 0x0201
		"00001010",	-- 0x0202
		"00000000",	-- 0x0203
		"01000011",	-- 0x0204
		"01101111",	-- 0x0205
		"01101100",	-- 0x0206
		"01100100",	-- 0x0207
		"00100000",	-- 0x0208
		"01110011",	-- 0x0209
		"01110100",	-- 0x020A
		"01100001",	-- 0x020B
		"01110010",	-- 0x020C
		"01110100",	-- 0x020D
		"00101100",	-- 0x020E
		"00100000",	-- 0x020F
		"01100011",	-- 0x0210
		"01101100",	-- 0x0211
		"01100101",	-- 0x0212
		"01100001",	-- 0x0213
		"01110010",	-- 0x0214
		"01101001",	-- 0x0215
		"01101110",	-- 0x0216
		"01100111",	-- 0x0217
		"00100000",	-- 0x0218
		"01101101",	-- 0x0219
		"01100101",	-- 0x021A
		"01101101",	-- 0x021B
		"01101111",	-- 0x021C
		"01110010",	-- 0x021D
		"01111001",	-- 0x021E
		"00101110",	-- 0x021F
		"00001101",	-- 0x0220
		"00001010",	-- 0x0221
		"00000000",	-- 0x0222
		"11001101",	-- 0x0223
		"11100001",	-- 0x0224
		"00001010",	-- 0x0225
		"11111110",	-- 0x0226
		"00001010",	-- 0x0227
		"00101000",	-- 0x0228
		"11111001",	-- 0x0229
		"11001101",	-- 0x022A
		"10111001",	-- 0x022B
		"00001010",	-- 0x022C
		"11111110",	-- 0x022D
		"00001101",	-- 0x022E
		"11000000",	-- 0x022F
		"00110011",	-- 0x0230
		"11000011",	-- 0x0231
		"01110100",	-- 0x0232
		"00000000",	-- 0x0233
		"11000101",	-- 0x0234
		"11010101",	-- 0x0235
		"11100101",	-- 0x0236
		"11111101",	-- 0x0237
		"11100101",	-- 0x0238
		"00100001",	-- 0x0239
		"01100001",	-- 0x023A
		"00000010",	-- 0x023B
		"11001101",	-- 0x023C
		"01101001",	-- 0x023D
		"00001011",	-- 0x023E
		"00100001",	-- 0x023F
		"01101101",	-- 0x0240
		"11111011",	-- 0x0241
		"00000110",	-- 0x0242
		"01010001",	-- 0x0243
		"11001101",	-- 0x0244
		"00010111",	-- 0x0245
		"00001011",	-- 0x0246
		"11111101",	-- 0x0247
		"00100001",	-- 0x0248
		"10111110",	-- 0x0249
		"11111011",	-- 0x024A
		"00010001",	-- 0x024B
		"01100001",	-- 0x024C
		"11111011",	-- 0x024D
		"11001101",	-- 0x024E
		"00110101",	-- 0x024F
		"00010000",	-- 0x0250
		"11001101",	-- 0x0251
		"01111010",	-- 0x0252
		"00001101",	-- 0x0253
		"00111000",	-- 0x0254
		"00000101",	-- 0x0255
		"11001101",	-- 0x0256
		"01100011",	-- 0x0257
		"00001011",	-- 0x0258
		"00011000",	-- 0x0259
		"11110110",	-- 0x025A
		"11111101",	-- 0x025B
		"11100001",	-- 0x025C
		"11100001",	-- 0x025D
		"11010001",	-- 0x025E
		"11000001",	-- 0x025F
		"11001001",	-- 0x0260
		"01000011",	-- 0x0261
		"01000001",	-- 0x0262
		"01010100",	-- 0x0263
		"00111010",	-- 0x0264
		"00100000",	-- 0x0265
		"01000110",	-- 0x0266
		"01001001",	-- 0x0267
		"01001100",	-- 0x0268
		"01000101",	-- 0x0269
		"01001110",	-- 0x026A
		"01000001",	-- 0x026B
		"01001101",	-- 0x026C
		"01000101",	-- 0x026D
		"00111101",	-- 0x026E
		"00000000",	-- 0x026F
		"11100101",	-- 0x0270
		"00100001",	-- 0x0271
		"01111100",	-- 0x0272
		"00000010",	-- 0x0273
		"11001101",	-- 0x0274
		"01101001",	-- 0x0275
		"00001011",	-- 0x0276
		"11001101",	-- 0x0277
		"10000110",	-- 0x0278
		"00010001",	-- 0x0279
		"11100001",	-- 0x027A
		"11001001",	-- 0x027B
		"01000100",	-- 0x027C
		"01001001",	-- 0x027D
		"01010010",	-- 0x027E
		"01000101",	-- 0x027F
		"01000011",	-- 0x0280
		"01010100",	-- 0x0281
		"01001111",	-- 0x0282
		"01010010",	-- 0x0283
		"01011001",	-- 0x0284
		"00001101",	-- 0x0285
		"00001010",	-- 0x0286
		"00000000",	-- 0x0287
		"11110101",	-- 0x0288
		"11100101",	-- 0x0289
		"00100001",	-- 0x028A
		"10101100",	-- 0x028B
		"00000010",	-- 0x028C
		"11001101",	-- 0x028D
		"01101001",	-- 0x028E
		"00001011",	-- 0x028F
		"11001101",	-- 0x0290
		"10001011",	-- 0x0291
		"00001011",	-- 0x0292
		"00100001",	-- 0x0293
		"00010011",	-- 0x0294
		"11111110",	-- 0x0295
		"00110110",	-- 0x0296
		"00001001",	-- 0x0297
		"11001101",	-- 0x0298
		"01101001",	-- 0x0299
		"00001011",	-- 0x029A
		"11001101",	-- 0x029B
		"11010100",	-- 0x029C
		"00001010",	-- 0x029D
		"00100001",	-- 0x029E
		"00101101",	-- 0x029F
		"11111110",	-- 0x02A0
		"00110110",	-- 0x02A1
		"00001001",	-- 0x02A2
		"11001101",	-- 0x02A3
		"01101001",	-- 0x02A4
		"00001011",	-- 0x02A5
		"11001101",	-- 0x02A6
		"11010100",	-- 0x02A7
		"00001010",	-- 0x02A8
		"11100001",	-- 0x02A9
		"11110001",	-- 0x02AA
		"11001001",	-- 0x02AB
		"01001001",	-- 0x02AC
		"01001110",	-- 0x02AD
		"01000110",	-- 0x02AE
		"01001111",	-- 0x02AF
		"00111010",	-- 0x02B0
		"00001101",	-- 0x02B1
		"00001010",	-- 0x02B2
		"00000000",	-- 0x02B3
		"11110101",	-- 0x02B4
		"11000101",	-- 0x02B5
		"11010101",	-- 0x02B6
		"11100101",	-- 0x02B7
		"11011101",	-- 0x02B8
		"11100101",	-- 0x02B9
		"00100001",	-- 0x02BA
		"00110011",	-- 0x02BB
		"00000011",	-- 0x02BC
		"11001101",	-- 0x02BD
		"01101001",	-- 0x02BE
		"00001011",	-- 0x02BF
		"11001101",	-- 0x02C0
		"11100001",	-- 0x02C1
		"00001010",	-- 0x02C2
		"11001101",	-- 0x02C3
		"10111001",	-- 0x02C4
		"00001010",	-- 0x02C5
		"11111110",	-- 0x02C6
		"01010010",	-- 0x02C7
		"00100000",	-- 0x02C8
		"00001001",	-- 0x02C9
		"11011101",	-- 0x02CA
		"00100001",	-- 0x02CB
		"00101011",	-- 0x02CC
		"00001100",	-- 0x02CD
		"00100001",	-- 0x02CE
		"00111101",	-- 0x02CF
		"00000011",	-- 0x02D0
		"00011000",	-- 0x02D1
		"00001011",	-- 0x02D2
		"11111110",	-- 0x02D3
		"01010111",	-- 0x02D4
		"00100000",	-- 0x02D5
		"11101001",	-- 0x02D6
		"11011101",	-- 0x02D7
		"00100001",	-- 0x02D8
		"10000010",	-- 0x02D9
		"00001100",	-- 0x02DA
		"00100001",	-- 0x02DB
		"01010111",	-- 0x02DC
		"00000011",	-- 0x02DD
		"11001101",	-- 0x02DE
		"01101001",	-- 0x02DF
		"00001011",	-- 0x02E0
		"11001101",	-- 0x02E1
		"00001100",	-- 0x02E2
		"00001011",	-- 0x02E3
		"11100101",	-- 0x02E4
		"00100001",	-- 0x02E5
		"01110010",	-- 0x02E6
		"00000011",	-- 0x02E7
		"11001101",	-- 0x02E8
		"01101001",	-- 0x02E9
		"00001011",	-- 0x02EA
		"11001101",	-- 0x02EB
		"11100111",	-- 0x02EC
		"00001010",	-- 0x02ED
		"11111110",	-- 0x02EE
		"00000000",	-- 0x02EF
		"00100000",	-- 0x02F0
		"00001000",	-- 0x02F1
		"00100001",	-- 0x02F2
		"10011111",	-- 0x02F3
		"00000011",	-- 0x02F4
		"11001101",	-- 0x02F5
		"01101001",	-- 0x02F6
		"00001011",	-- 0x02F7
		"00011000",	-- 0x02F8
		"00110000",	-- 0x02F9
		"00100001",	-- 0x02FA
		"10010000",	-- 0x02FB
		"00000011",	-- 0x02FC
		"11001101",	-- 0x02FD
		"01101001",	-- 0x02FE
		"00001011",	-- 0x02FF
		"11001101",	-- 0x0300
		"00001100",	-- 0x0301
		"00001011",	-- 0x0302
		"01000100",	-- 0x0303
		"01001101",	-- 0x0304
		"11001101",	-- 0x0305
		"00001100",	-- 0x0306
		"00001011",	-- 0x0307
		"01010100",	-- 0x0308
		"01011101",	-- 0x0309
		"11100001",	-- 0x030A
		"11110101",	-- 0x030B
		"11001101",	-- 0x030C
		"00110001",	-- 0x030D
		"00000011",	-- 0x030E
		"11100101",	-- 0x030F
		"11000101",	-- 0x0310
		"01100010",	-- 0x0311
		"01101011",	-- 0x0312
		"00000001",	-- 0x0313
		"00000001",	-- 0x0314
		"00000000",	-- 0x0315
		"00001001",	-- 0x0316
		"01010100",	-- 0x0317
		"01011101",	-- 0x0318
		"11100001",	-- 0x0319
		"00110000",	-- 0x031A
		"00000001",	-- 0x031B
		"00001001",	-- 0x031C
		"01000100",	-- 0x031D
		"01001101",	-- 0x031E
		"11100001",	-- 0x031F
		"11000101",	-- 0x0320
		"00000001",	-- 0x0321
		"00000000",	-- 0x0322
		"00000010",	-- 0x0323
		"00001001",	-- 0x0324
		"11000001",	-- 0x0325
		"11110001",	-- 0x0326
		"00111101",	-- 0x0327
		"00100000",	-- 0x0328
		"11100001",	-- 0x0329
		"11011101",	-- 0x032A
		"11100001",	-- 0x032B
		"11100001",	-- 0x032C
		"11010001",	-- 0x032D
		"11000001",	-- 0x032E
		"11110001",	-- 0x032F
		"11001001",	-- 0x0330
		"11011101",	-- 0x0331
		"11101001",	-- 0x0332
		"01010100",	-- 0x0333
		"01010010",	-- 0x0334
		"01000001",	-- 0x0335
		"01001110",	-- 0x0336
		"01010011",	-- 0x0337
		"01000110",	-- 0x0338
		"01000101",	-- 0x0339
		"01010010",	-- 0x033A
		"00101111",	-- 0x033B
		"00000000",	-- 0x033C
		"01010010",	-- 0x033D
		"01000101",	-- 0x033E
		"01000001",	-- 0x033F
		"01000100",	-- 0x0340
		"00111010",	-- 0x0341
		"00100000",	-- 0x0342
		"00001101",	-- 0x0343
		"00001010",	-- 0x0344
		"00100000",	-- 0x0345
		"00100000",	-- 0x0346
		"00100000",	-- 0x0347
		"00100000",	-- 0x0348
		"01001101",	-- 0x0349
		"01000101",	-- 0x034A
		"01001101",	-- 0x034B
		"01001111",	-- 0x034C
		"01010010",	-- 0x034D
		"01011001",	-- 0x034E
		"00100000",	-- 0x034F
		"01010011",	-- 0x0350
		"01010100",	-- 0x0351
		"01000001",	-- 0x0352
		"01010010",	-- 0x0353
		"01010100",	-- 0x0354
		"00111101",	-- 0x0355
		"00000000",	-- 0x0356
		"01010111",	-- 0x0357
		"01010010",	-- 0x0358
		"01001001",	-- 0x0359
		"01010100",	-- 0x035A
		"01000101",	-- 0x035B
		"00111010",	-- 0x035C
		"00100000",	-- 0x035D
		"00001101",	-- 0x035E
		"00001010",	-- 0x035F
		"00100000",	-- 0x0360
		"00100000",	-- 0x0361
		"00100000",	-- 0x0362
		"00100000",	-- 0x0363
		"01001101",	-- 0x0364
		"01000101",	-- 0x0365
		"01001101",	-- 0x0366
		"01001111",	-- 0x0367
		"01010010",	-- 0x0368
		"01011001",	-- 0x0369
		"00100000",	-- 0x036A
		"01010011",	-- 0x036B
		"01010100",	-- 0x036C
		"01000001",	-- 0x036D
		"01010010",	-- 0x036E
		"01010100",	-- 0x036F
		"00111101",	-- 0x0370
		"00000000",	-- 0x0371
		"00100000",	-- 0x0372
		"01001110",	-- 0x0373
		"01010101",	-- 0x0374
		"01001101",	-- 0x0375
		"01000010",	-- 0x0376
		"01000101",	-- 0x0377
		"01010010",	-- 0x0378
		"00100000",	-- 0x0379
		"01001111",	-- 0x037A
		"01000110",	-- 0x037B
		"00100000",	-- 0x037C
		"01000010",	-- 0x037D
		"01001100",	-- 0x037E
		"01001111",	-- 0x037F
		"01000011",	-- 0x0380
		"01001011",	-- 0x0381
		"01010011",	-- 0x0382
		"00100000",	-- 0x0383
		"00101000",	-- 0x0384
		"00110101",	-- 0x0385
		"00110001",	-- 0x0386
		"00110010",	-- 0x0387
		"00100000",	-- 0x0388
		"01000010",	-- 0x0389
		"01011001",	-- 0x038A
		"01010100",	-- 0x038B
		"01000101",	-- 0x038C
		"00101001",	-- 0x038D
		"00111101",	-- 0x038E
		"00000000",	-- 0x038F
		"00100000",	-- 0x0390
		"01010011",	-- 0x0391
		"01010100",	-- 0x0392
		"01000001",	-- 0x0393
		"01010010",	-- 0x0394
		"01010100",	-- 0x0395
		"00100000",	-- 0x0396
		"01010011",	-- 0x0397
		"01000101",	-- 0x0398
		"01000011",	-- 0x0399
		"01010100",	-- 0x039A
		"01001111",	-- 0x039B
		"01010010",	-- 0x039C
		"00111101",	-- 0x039D
		"00000000",	-- 0x039E
		"00100000",	-- 0x039F
		"01001110",	-- 0x03A0
		"01101111",	-- 0x03A1
		"01110100",	-- 0x03A2
		"01101000",	-- 0x03A3
		"01101001",	-- 0x03A4
		"01101110",	-- 0x03A5
		"01100111",	-- 0x03A6
		"00100000",	-- 0x03A7
		"01110100",	-- 0x03A8
		"01101111",	-- 0x03A9
		"00100000",	-- 0x03AA
		"01100100",	-- 0x03AB
		"01101111",	-- 0x03AC
		"00100000",	-- 0x03AD
		"01100110",	-- 0x03AE
		"01101111",	-- 0x03AF
		"01110010",	-- 0x03B0
		"00100000",	-- 0x03B1
		"01111010",	-- 0x03B2
		"01100101",	-- 0x03B3
		"01110010",	-- 0x03B4
		"01101111",	-- 0x03B5
		"00100000",	-- 0x03B6
		"01100010",	-- 0x03B7
		"01101100",	-- 0x03B8
		"01101111",	-- 0x03B9
		"01100011",	-- 0x03BA
		"01101011",	-- 0x03BB
		"01110011",	-- 0x03BC
		"00101110",	-- 0x03BD
		"00001101",	-- 0x03BE
		"00001010",	-- 0x03BF
		"00000000",	-- 0x03C0
		"11110101",	-- 0x03C1
		"11000101",	-- 0x03C2
		"11010101",	-- 0x03C3
		"11100101",	-- 0x03C4
		"00100001",	-- 0x03C5
		"00100001",	-- 0x03C6
		"00000100",	-- 0x03C7
		"11001101",	-- 0x03C8
		"01101001",	-- 0x03C9
		"00001011",	-- 0x03CA
		"11001101",	-- 0x03CB
		"00001100",	-- 0x03CC
		"00001011",	-- 0x03CD
		"11100101",	-- 0x03CE
		"00100001",	-- 0x03CF
		"00101110",	-- 0x03D0
		"00000100",	-- 0x03D1
		"11001101",	-- 0x03D2
		"01101001",	-- 0x03D3
		"00001011",	-- 0x03D4
		"11001101",	-- 0x03D5
		"00001100",	-- 0x03D6
		"00001011",	-- 0x03D7
		"11001101",	-- 0x03D8
		"11010100",	-- 0x03D9
		"00001010",	-- 0x03DA
		"00100011",	-- 0x03DB
		"01010100",	-- 0x03DC
		"01011101",	-- 0x03DD
		"11100001",	-- 0x03DE
		"00000110",	-- 0x03DF
		"00010000",	-- 0x03E0
		"11100101",	-- 0x03E1
		"11001101",	-- 0x03E2
		"01010110",	-- 0x03E3
		"00001011",	-- 0x03E4
		"00100001",	-- 0x03E5
		"00110100",	-- 0x03E6
		"00000100",	-- 0x03E7
		"11001101",	-- 0x03E8
		"01101001",	-- 0x03E9
		"00001011",	-- 0x03EA
		"11100001",	-- 0x03EB
		"11100101",	-- 0x03EC
		"01111110",	-- 0x03ED
		"11001101",	-- 0x03EE
		"00110101",	-- 0x03EF
		"00001011",	-- 0x03F0
		"00111110",	-- 0x03F1
		"00100000",	-- 0x03F2
		"11001101",	-- 0x03F3
		"01100011",	-- 0x03F4
		"00001011",	-- 0x03F5
		"00100011",	-- 0x03F6
		"00010000",	-- 0x03F7
		"11110100",	-- 0x03F8
		"00000110",	-- 0x03F9
		"00010000",	-- 0x03FA
		"00111110",	-- 0x03FB
		"00100000",	-- 0x03FC
		"11001101",	-- 0x03FD
		"01100011",	-- 0x03FE
		"00001011",	-- 0x03FF
		"11001101",	-- 0x0400
		"01100011",	-- 0x0401
		"00001011",	-- 0x0402
		"11100001",	-- 0x0403
		"01111110",	-- 0x0404
		"11001101",	-- 0x0405
		"10100101",	-- 0x0406
		"00001010",	-- 0x0407
		"00111000",	-- 0x0408
		"00000010",	-- 0x0409
		"00111110",	-- 0x040A
		"00101110",	-- 0x040B
		"11001101",	-- 0x040C
		"01100011",	-- 0x040D
		"00001011",	-- 0x040E
		"00100011",	-- 0x040F
		"00010000",	-- 0x0410
		"11110010",	-- 0x0411
		"11001101",	-- 0x0412
		"11010100",	-- 0x0413
		"00001010",	-- 0x0414
		"11100101",	-- 0x0415
		"10100111",	-- 0x0416
		"11101101",	-- 0x0417
		"01010010",	-- 0x0418
		"11100001",	-- 0x0419
		"00111000",	-- 0x041A
		"11000011",	-- 0x041B
		"11100001",	-- 0x041C
		"11010001",	-- 0x041D
		"11000001",	-- 0x041E
		"11110001",	-- 0x041F
		"11001001",	-- 0x0420
		"01000100",	-- 0x0421
		"01010101",	-- 0x0422
		"01001101",	-- 0x0423
		"01010000",	-- 0x0424
		"00111010",	-- 0x0425
		"00100000",	-- 0x0426
		"01010011",	-- 0x0427
		"01010100",	-- 0x0428
		"01000001",	-- 0x0429
		"01010010",	-- 0x042A
		"01010100",	-- 0x042B
		"00111101",	-- 0x042C
		"00000000",	-- 0x042D
		"00100000",	-- 0x042E
		"01000101",	-- 0x042F
		"01001110",	-- 0x0430
		"01000100",	-- 0x0431
		"00111101",	-- 0x0432
		"00000000",	-- 0x0433
		"00111010",	-- 0x0434
		"00100000",	-- 0x0435
		"00000000",	-- 0x0436
		"11110101",	-- 0x0437
		"11100101",	-- 0x0438
		"00100001",	-- 0x0439
		"01100101",	-- 0x043A
		"00000100",	-- 0x043B
		"11001101",	-- 0x043C
		"01101001",	-- 0x043D
		"00001011",	-- 0x043E
		"11001101",	-- 0x043F
		"00001100",	-- 0x0440
		"00001011",	-- 0x0441
		"11100101",	-- 0x0442
		"00100001",	-- 0x0443
		"10000011",	-- 0x0444
		"00000100",	-- 0x0445
		"11001101",	-- 0x0446
		"01101001",	-- 0x0447
		"00001011",	-- 0x0448
		"11100001",	-- 0x0449
		"01111110",	-- 0x044A
		"00100011",	-- 0x044B
		"11100101",	-- 0x044C
		"11001101",	-- 0x044D
		"00110101",	-- 0x044E
		"00001011",	-- 0x044F
		"11001101",	-- 0x0450
		"11100001",	-- 0x0451
		"00001010",	-- 0x0452
		"11111110",	-- 0x0453
		"00100000",	-- 0x0454
		"00100000",	-- 0x0455
		"00000111",	-- 0x0456
		"00111110",	-- 0x0457
		"00100000",	-- 0x0458
		"11001101",	-- 0x0459
		"01100011",	-- 0x045A
		"00001011",	-- 0x045B
		"00011000",	-- 0x045C
		"11101011",	-- 0x045D
		"11100001",	-- 0x045E
		"11001101",	-- 0x045F
		"11010100",	-- 0x0460
		"00001010",	-- 0x0461
		"11100001",	-- 0x0462
		"11110001",	-- 0x0463
		"11001001",	-- 0x0464
		"01000101",	-- 0x0465
		"01011000",	-- 0x0466
		"01000001",	-- 0x0467
		"01001101",	-- 0x0468
		"01001001",	-- 0x0469
		"01001110",	-- 0x046A
		"01000101",	-- 0x046B
		"00100000",	-- 0x046C
		"00101000",	-- 0x046D
		"01110100",	-- 0x046E
		"01111001",	-- 0x046F
		"01110000",	-- 0x0470
		"01100101",	-- 0x0471
		"00100000",	-- 0x0472
		"00100111",	-- 0x0473
		"00100000",	-- 0x0474
		"00100111",	-- 0x0475
		"00101111",	-- 0x0476
		"01010010",	-- 0x0477
		"01000101",	-- 0x0478
		"01010100",	-- 0x0479
		"00101001",	-- 0x047A
		"00111010",	-- 0x047B
		"00100000",	-- 0x047C
		"01000001",	-- 0x047D
		"01000100",	-- 0x047E
		"01000100",	-- 0x047F
		"01010010",	-- 0x0480
		"00111101",	-- 0x0481
		"00000000",	-- 0x0482
		"00100000",	-- 0x0483
		"01000100",	-- 0x0484
		"01000001",	-- 0x0485
		"01010100",	-- 0x0486
		"01000001",	-- 0x0487
		"00111101",	-- 0x0488
		"00000000",	-- 0x0489
		"11110101",	-- 0x048A
		"11000101",	-- 0x048B
		"11010101",	-- 0x048C
		"11100101",	-- 0x048D
		"00100001",	-- 0x048E
		"11100100",	-- 0x048F
		"00000100",	-- 0x0490
		"11001101",	-- 0x0491
		"01101001",	-- 0x0492
		"00001011",	-- 0x0493
		"11001101",	-- 0x0494
		"00001100",	-- 0x0495
		"00001011",	-- 0x0496
		"11100101",	-- 0x0497
		"10100111",	-- 0x0498
		"00000001",	-- 0x0499
		"00000000",	-- 0x049A
		"10000000",	-- 0x049B
		"11101101",	-- 0x049C
		"01000010",	-- 0x049D
		"00110000",	-- 0x049E
		"00001001",	-- 0x049F
		"00100001",	-- 0x04A0
		"00000010",	-- 0x04A1
		"00000101",	-- 0x04A2
		"11001101",	-- 0x04A3
		"01101001",	-- 0x04A4
		"00001011",	-- 0x04A5
		"11100001",	-- 0x04A6
		"00011000",	-- 0x04A7
		"00110110",	-- 0x04A8
		"00100001",	-- 0x04A9
		"11110001",	-- 0x04AA
		"00000100",	-- 0x04AB
		"11001101",	-- 0x04AC
		"01101001",	-- 0x04AD
		"00001011",	-- 0x04AE
		"11001101",	-- 0x04AF
		"00001100",	-- 0x04B0
		"00001011",	-- 0x04B1
		"01000100",	-- 0x04B2
		"01001101",	-- 0x04B3
		"11100001",	-- 0x04B4
		"11100101",	-- 0x04B5
		"11000101",	-- 0x04B6
		"00001001",	-- 0x04B7
		"10100111",	-- 0x04B8
		"00000001",	-- 0x04B9
		"00000000",	-- 0x04BA
		"10000000",	-- 0x04BB
		"11101101",	-- 0x04BC
		"01000010",	-- 0x04BD
		"00110000",	-- 0x04BE
		"00001010",	-- 0x04BF
		"00100001",	-- 0x04C0
		"00010110",	-- 0x04C1
		"00000101",	-- 0x04C2
		"11001101",	-- 0x04C3
		"01101001",	-- 0x04C4
		"00001011",	-- 0x04C5
		"11000001",	-- 0x04C6
		"11100001",	-- 0x04C7
		"00011000",	-- 0x04C8
		"00010101",	-- 0x04C9
		"00100001",	-- 0x04CA
		"11111010",	-- 0x04CB
		"00000100",	-- 0x04CC
		"11001101",	-- 0x04CD
		"01101001",	-- 0x04CE
		"00001011",	-- 0x04CF
		"11001101",	-- 0x04D0
		"11100111",	-- 0x04D1
		"00001010",	-- 0x04D2
		"11000001",	-- 0x04D3
		"11100001",	-- 0x04D4
		"01010100",	-- 0x04D5
		"01011101",	-- 0x04D6
		"00010011",	-- 0x04D7
		"00001011",	-- 0x04D8
		"01110111",	-- 0x04D9
		"11101101",	-- 0x04DA
		"10110000",	-- 0x04DB
		"11001101",	-- 0x04DC
		"11010100",	-- 0x04DD
		"00001010",	-- 0x04DE
		"11100001",	-- 0x04DF
		"11010001",	-- 0x04E0
		"11000001",	-- 0x04E1
		"11110001",	-- 0x04E2
		"11001001",	-- 0x04E3
		"01000110",	-- 0x04E4
		"01001001",	-- 0x04E5
		"01001100",	-- 0x04E6
		"01001100",	-- 0x04E7
		"00111010",	-- 0x04E8
		"00100000",	-- 0x04E9
		"01010011",	-- 0x04EA
		"01010100",	-- 0x04EB
		"01000001",	-- 0x04EC
		"01010010",	-- 0x04ED
		"01010100",	-- 0x04EE
		"00111101",	-- 0x04EF
		"00000000",	-- 0x04F0
		"00100000",	-- 0x04F1
		"01001100",	-- 0x04F2
		"01000101",	-- 0x04F3
		"01001110",	-- 0x04F4
		"01000111",	-- 0x04F5
		"01010100",	-- 0x04F6
		"01001000",	-- 0x04F7
		"00111101",	-- 0x04F8
		"00000000",	-- 0x04F9
		"00100000",	-- 0x04FA
		"01010110",	-- 0x04FB
		"01000001",	-- 0x04FC
		"01001100",	-- 0x04FD
		"01010101",	-- 0x04FE
		"01000101",	-- 0x04FF
		"00111101",	-- 0x0500
		"00000000",	-- 0x0501
		"00100000",	-- 0x0502
		"01001001",	-- 0x0503
		"01101100",	-- 0x0504
		"01101100",	-- 0x0505
		"01100101",	-- 0x0506
		"01100111",	-- 0x0507
		"01100001",	-- 0x0508
		"01101100",	-- 0x0509
		"00100000",	-- 0x050A
		"01100001",	-- 0x050B
		"01100100",	-- 0x050C
		"01100100",	-- 0x050D
		"01110010",	-- 0x050E
		"01100101",	-- 0x050F
		"01110011",	-- 0x0510
		"01110011",	-- 0x0511
		"00100001",	-- 0x0512
		"00001101",	-- 0x0513
		"00001010",	-- 0x0514
		"00000000",	-- 0x0515
		"00100000",	-- 0x0516
		"01000010",	-- 0x0517
		"01101100",	-- 0x0518
		"01101111",	-- 0x0519
		"01100011",	-- 0x051A
		"01101011",	-- 0x051B
		"00100000",	-- 0x051C
		"01100101",	-- 0x051D
		"01111000",	-- 0x051E
		"01100011",	-- 0x051F
		"01100101",	-- 0x0520
		"01100101",	-- 0x0521
		"01100100",	-- 0x0522
		"01110011",	-- 0x0523
		"00100000",	-- 0x0524
		"01010010",	-- 0x0525
		"01000001",	-- 0x0526
		"01001101",	-- 0x0527
		"00100000",	-- 0x0528
		"01100001",	-- 0x0529
		"01110010",	-- 0x052A
		"01100101",	-- 0x052B
		"01100001",	-- 0x052C
		"00100001",	-- 0x052D
		"00001101",	-- 0x052E
		"00001010",	-- 0x052F
		"00000000",	-- 0x0530
		"11100101",	-- 0x0531
		"00100001",	-- 0x0532
		"00111010",	-- 0x0533
		"00000101",	-- 0x0534
		"11001101",	-- 0x0535
		"01101001",	-- 0x0536
		"00001011",	-- 0x0537
		"11100001",	-- 0x0538
		"11001001",	-- 0x0539
		"01001000",	-- 0x053A
		"01000101",	-- 0x053B
		"01001100",	-- 0x053C
		"01010000",	-- 0x053D
		"00111010",	-- 0x053E
		"00100000",	-- 0x053F
		"01001011",	-- 0x0540
		"01101110",	-- 0x0541
		"01101111",	-- 0x0542
		"01110111",	-- 0x0543
		"01101110",	-- 0x0544
		"00100000",	-- 0x0545
		"01100011",	-- 0x0546
		"01101111",	-- 0x0547
		"01101101",	-- 0x0548
		"01101101",	-- 0x0549
		"01100001",	-- 0x054A
		"01101110",	-- 0x054B
		"01100100",	-- 0x054C
		"00100000",	-- 0x054D
		"01100111",	-- 0x054E
		"01110010",	-- 0x054F
		"01101111",	-- 0x0550
		"01110101",	-- 0x0551
		"01110000",	-- 0x0552
		"01110011",	-- 0x0553
		"00100000",	-- 0x0554
		"01100001",	-- 0x0555
		"01101110",	-- 0x0556
		"01100100",	-- 0x0557
		"00100000",	-- 0x0558
		"01100011",	-- 0x0559
		"01101111",	-- 0x055A
		"01101101",	-- 0x055B
		"01101101",	-- 0x055C
		"01100001",	-- 0x055D
		"01101110",	-- 0x055E
		"01100100",	-- 0x055F
		"01110011",	-- 0x0560
		"00111010",	-- 0x0561
		"00001101",	-- 0x0562
		"00001010",	-- 0x0563
		"00100000",	-- 0x0564
		"00100000",	-- 0x0565
		"00100000",	-- 0x0566
		"00100000",	-- 0x0567
		"00100000",	-- 0x0568
		"00100000",	-- 0x0569
		"00100000",	-- 0x056A
		"00100000",	-- 0x056B
		"00100000",	-- 0x056C
		"01000011",	-- 0x056D
		"00101000",	-- 0x056E
		"01101111",	-- 0x056F
		"01101110",	-- 0x0570
		"01110100",	-- 0x0571
		"01110010",	-- 0x0572
		"01101111",	-- 0x0573
		"01101100",	-- 0x0574
		"00100000",	-- 0x0575
		"01100111",	-- 0x0576
		"01110010",	-- 0x0577
		"01101111",	-- 0x0578
		"01110101",	-- 0x0579
		"01110000",	-- 0x057A
		"00101001",	-- 0x057B
		"00111010",	-- 0x057C
		"00001101",	-- 0x057D
		"00001010",	-- 0x057E
		"00100000",	-- 0x057F
		"00100000",	-- 0x0580
		"00100000",	-- 0x0581
		"00100000",	-- 0x0582
		"00100000",	-- 0x0583
		"00100000",	-- 0x0584
		"00100000",	-- 0x0585
		"00100000",	-- 0x0586
		"00100000",	-- 0x0587
		"00100000",	-- 0x0588
		"00100000",	-- 0x0589
		"00100000",	-- 0x058A
		"00100000",	-- 0x058B
		"01000011",	-- 0x058C
		"00101000",	-- 0x058D
		"01101111",	-- 0x058E
		"01101100",	-- 0x058F
		"01100100",	-- 0x0590
		"00100000",	-- 0x0591
		"01110011",	-- 0x0592
		"01110100",	-- 0x0593
		"01100001",	-- 0x0594
		"01110010",	-- 0x0595
		"01110100",	-- 0x0596
		"00101001",	-- 0x0597
		"00101100",	-- 0x0598
		"00100000",	-- 0x0599
		"01001001",	-- 0x059A
		"00101000",	-- 0x059B
		"01101110",	-- 0x059C
		"01100110",	-- 0x059D
		"01101111",	-- 0x059E
		"00101001",	-- 0x059F
		"00101100",	-- 0x05A0
		"00100000",	-- 0x05A1
		"01010011",	-- 0x05A2
		"00101000",	-- 0x05A3
		"01110100",	-- 0x05A4
		"01100001",	-- 0x05A5
		"01110010",	-- 0x05A6
		"01110100",	-- 0x05A7
		"00101001",	-- 0x05A8
		"00101100",	-- 0x05A9
		"00100000",	-- 0x05AA
		"01010111",	-- 0x05AB
		"00101000",	-- 0x05AC
		"01100001",	-- 0x05AD
		"01110010",	-- 0x05AE
		"01101101",	-- 0x05AF
		"00100000",	-- 0x05B0
		"01110011",	-- 0x05B1
		"01110100",	-- 0x05B2
		"01100001",	-- 0x05B3
		"01110010",	-- 0x05B4
		"01110100",	-- 0x05B5
		"00101001",	-- 0x05B6
		"00001101",	-- 0x05B7
		"00001010",	-- 0x05B8
		"00100000",	-- 0x05B9
		"00100000",	-- 0x05BA
		"00100000",	-- 0x05BB
		"00100000",	-- 0x05BC
		"00100000",	-- 0x05BD
		"00100000",	-- 0x05BE
		"00100000",	-- 0x05BF
		"00100000",	-- 0x05C0
		"00100000",	-- 0x05C1
		"01000100",	-- 0x05C2
		"00101000",	-- 0x05C3
		"01101001",	-- 0x05C4
		"01110011",	-- 0x05C5
		"01101011",	-- 0x05C6
		"00100000",	-- 0x05C7
		"01100111",	-- 0x05C8
		"01110010",	-- 0x05C9
		"01101111",	-- 0x05CA
		"01110101",	-- 0x05CB
		"01110000",	-- 0x05CC
		"00101001",	-- 0x05CD
		"00111010",	-- 0x05CE
		"00001101",	-- 0x05CF
		"00001010",	-- 0x05D0
		"00100000",	-- 0x05D1
		"00100000",	-- 0x05D2
		"00100000",	-- 0x05D3
		"00100000",	-- 0x05D4
		"00100000",	-- 0x05D5
		"00100000",	-- 0x05D6
		"00100000",	-- 0x05D7
		"00100000",	-- 0x05D8
		"00100000",	-- 0x05D9
		"00100000",	-- 0x05DA
		"00100000",	-- 0x05DB
		"00100000",	-- 0x05DC
		"00100000",	-- 0x05DD
		"01001001",	-- 0x05DE
		"00101000",	-- 0x05DF
		"01101110",	-- 0x05E0
		"01100110",	-- 0x05E1
		"01101111",	-- 0x05E2
		"00101001",	-- 0x05E3
		"00101100",	-- 0x05E4
		"00100000",	-- 0x05E5
		"01001101",	-- 0x05E6
		"00101000",	-- 0x05E7
		"01101111",	-- 0x05E8
		"01110101",	-- 0x05E9
		"01101110",	-- 0x05EA
		"01110100",	-- 0x05EB
		"00101001",	-- 0x05EC
		"00101100",	-- 0x05ED
		"00100000",	-- 0x05EE
		"01010100",	-- 0x05EF
		"00101000",	-- 0x05F0
		"01110010",	-- 0x05F1
		"01100001",	-- 0x05F2
		"01101110",	-- 0x05F3
		"01110011",	-- 0x05F4
		"01100110",	-- 0x05F5
		"01100101",	-- 0x05F6
		"01110010",	-- 0x05F7
		"00101001",	-- 0x05F8
		"00101100",	-- 0x05F9
		"00100000",	-- 0x05FA
		"00100000",	-- 0x05FB
		"00100000",	-- 0x05FC
		"00100000",	-- 0x05FD
		"00100000",	-- 0x05FE
		"00100000",	-- 0x05FF
		"00100000",	-- 0x0600
		"00100000",	-- 0x0601
		"00100000",	-- 0x0602
		"01010101",	-- 0x0603
		"00101000",	-- 0x0604
		"01101110",	-- 0x0605
		"01101101",	-- 0x0606
		"01101111",	-- 0x0607
		"01110101",	-- 0x0608
		"01101110",	-- 0x0609
		"01110100",	-- 0x060A
		"00101001",	-- 0x060B
		"00001101",	-- 0x060C
		"00001010",	-- 0x060D
		"00100000",	-- 0x060E
		"00100000",	-- 0x060F
		"00100000",	-- 0x0610
		"00100000",	-- 0x0611
		"00100000",	-- 0x0612
		"00100000",	-- 0x0613
		"00100000",	-- 0x0614
		"00100000",	-- 0x0615
		"00100000",	-- 0x0616
		"00100000",	-- 0x0617
		"00100000",	-- 0x0618
		"00100000",	-- 0x0619
		"00100000",	-- 0x061A
		"00100000",	-- 0x061B
		"00100000",	-- 0x061C
		"00100000",	-- 0x061D
		"00100000",	-- 0x061E
		"00100000",	-- 0x061F
		"00100000",	-- 0x0620
		"00100000",	-- 0x0621
		"00100000",	-- 0x0622
		"00100000",	-- 0x0623
		"00100000",	-- 0x0624
		"00100000",	-- 0x0625
		"00100000",	-- 0x0626
		"00100000",	-- 0x0627
		"00100000",	-- 0x0628
		"00100000",	-- 0x0629
		"00100000",	-- 0x062A
		"00100000",	-- 0x062B
		"00100000",	-- 0x062C
		"00100000",	-- 0x062D
		"00100000",	-- 0x062E
		"00100000",	-- 0x062F
		"01010010",	-- 0x0630
		"00101000",	-- 0x0631
		"01100101",	-- 0x0632
		"01100001",	-- 0x0633
		"01100100",	-- 0x0634
		"00101001",	-- 0x0635
		"00101100",	-- 0x0636
		"00100000",	-- 0x0637
		"01010111",	-- 0x0638
		"00101000",	-- 0x0639
		"01110010",	-- 0x063A
		"01101001",	-- 0x063B
		"01110100",	-- 0x063C
		"01100101",	-- 0x063D
		"00101001",	-- 0x063E
		"00001101",	-- 0x063F
		"00001010",	-- 0x0640
		"00100000",	-- 0x0641
		"00100000",	-- 0x0642
		"00100000",	-- 0x0643
		"00100000",	-- 0x0644
		"00100000",	-- 0x0645
		"00100000",	-- 0x0646
		"00100000",	-- 0x0647
		"00100000",	-- 0x0648
		"00100000",	-- 0x0649
		"01000110",	-- 0x064A
		"00101000",	-- 0x064B
		"01101001",	-- 0x064C
		"01101100",	-- 0x064D
		"01100101",	-- 0x064E
		"00100000",	-- 0x064F
		"01100111",	-- 0x0650
		"01110010",	-- 0x0651
		"01101111",	-- 0x0652
		"01110101",	-- 0x0653
		"01110000",	-- 0x0654
		"00101001",	-- 0x0655
		"00111010",	-- 0x0656
		"00001101",	-- 0x0657
		"00001010",	-- 0x0658
		"00100000",	-- 0x0659
		"00100000",	-- 0x065A
		"00100000",	-- 0x065B
		"00100000",	-- 0x065C
		"00100000",	-- 0x065D
		"00100000",	-- 0x065E
		"00100000",	-- 0x065F
		"00100000",	-- 0x0660
		"00100000",	-- 0x0661
		"00100000",	-- 0x0662
		"00100000",	-- 0x0663
		"00100000",	-- 0x0664
		"00100000",	-- 0x0665
		"01000011",	-- 0x0666
		"00101000",	-- 0x0667
		"01100001",	-- 0x0668
		"01110100",	-- 0x0669
		"00101001",	-- 0x066A
		"00101100",	-- 0x066B
		"00100000",	-- 0x066C
		"01000100",	-- 0x066D
		"00101000",	-- 0x066E
		"01101001",	-- 0x066F
		"01110010",	-- 0x0670
		"01100101",	-- 0x0671
		"01100011",	-- 0x0672
		"01110100",	-- 0x0673
		"01101111",	-- 0x0674
		"01110010",	-- 0x0675
		"01111001",	-- 0x0676
		"00101001",	-- 0x0677
		"00101100",	-- 0x0678
		"00100000",	-- 0x0679
		"01001100",	-- 0x067A
		"00101000",	-- 0x067B
		"01101111",	-- 0x067C
		"01100001",	-- 0x067D
		"01100100",	-- 0x067E
		"00101001",	-- 0x067F
		"00001101",	-- 0x0680
		"00001010",	-- 0x0681
		"00100000",	-- 0x0682
		"00100000",	-- 0x0683
		"00100000",	-- 0x0684
		"00100000",	-- 0x0685
		"00100000",	-- 0x0686
		"00100000",	-- 0x0687
		"00100000",	-- 0x0688
		"00100000",	-- 0x0689
		"00100000",	-- 0x068A
		"01001000",	-- 0x068B
		"00101000",	-- 0x068C
		"01100101",	-- 0x068D
		"01101100",	-- 0x068E
		"01110000",	-- 0x068F
		"00101001",	-- 0x0690
		"00001101",	-- 0x0691
		"00001010",	-- 0x0692
		"00100000",	-- 0x0693
		"00100000",	-- 0x0694
		"00100000",	-- 0x0695
		"00100000",	-- 0x0696
		"00100000",	-- 0x0697
		"00100000",	-- 0x0698
		"00100000",	-- 0x0699
		"00100000",	-- 0x069A
		"00100000",	-- 0x069B
		"01001101",	-- 0x069C
		"00101000",	-- 0x069D
		"01100101",	-- 0x069E
		"01101101",	-- 0x069F
		"01101111",	-- 0x06A0
		"01110010",	-- 0x06A1
		"01111001",	-- 0x06A2
		"00100000",	-- 0x06A3
		"01100111",	-- 0x06A4
		"01110010",	-- 0x06A5
		"01101111",	-- 0x06A6
		"01110101",	-- 0x06A7
		"01110000",	-- 0x06A8
		"00101001",	-- 0x06A9
		"00111010",	-- 0x06AA
		"00001101",	-- 0x06AB
		"00001010",	-- 0x06AC
		"00100000",	-- 0x06AD
		"00100000",	-- 0x06AE
		"00100000",	-- 0x06AF
		"00100000",	-- 0x06B0
		"00100000",	-- 0x06B1
		"00100000",	-- 0x06B2
		"00100000",	-- 0x06B3
		"00100000",	-- 0x06B4
		"00100000",	-- 0x06B5
		"00100000",	-- 0x06B6
		"00100000",	-- 0x06B7
		"00100000",	-- 0x06B8
		"00100000",	-- 0x06B9
		"01000100",	-- 0x06BA
		"00101000",	-- 0x06BB
		"01110101",	-- 0x06BC
		"01101101",	-- 0x06BD
		"01110000",	-- 0x06BE
		"00101001",	-- 0x06BF
		"00101100",	-- 0x06C0
		"00100000",	-- 0x06C1
		"01000101",	-- 0x06C2
		"00101000",	-- 0x06C3
		"01111000",	-- 0x06C4
		"01100001",	-- 0x06C5
		"01101101",	-- 0x06C6
		"01101001",	-- 0x06C7
		"01101110",	-- 0x06C8
		"01100101",	-- 0x06C9
		"00101001",	-- 0x06CA
		"00101100",	-- 0x06CB
		"00100000",	-- 0x06CC
		"01000110",	-- 0x06CD
		"00101000",	-- 0x06CE
		"01101001",	-- 0x06CF
		"01101100",	-- 0x06D0
		"01101100",	-- 0x06D1
		"00101001",	-- 0x06D2
		"00101100",	-- 0x06D3
		"00100000",	-- 0x06D4
		"01001001",	-- 0x06D5
		"00101000",	-- 0x06D6
		"01101110",	-- 0x06D7
		"01110100",	-- 0x06D8
		"01100101",	-- 0x06D9
		"01101100",	-- 0x06DA
		"00100000",	-- 0x06DB
		"01001000",	-- 0x06DC
		"01100101",	-- 0x06DD
		"01111000",	-- 0x06DE
		"00100000",	-- 0x06DF
		"01001100",	-- 0x06E0
		"01101111",	-- 0x06E1
		"01100001",	-- 0x06E2
		"01100100",	-- 0x06E3
		"00101001",	-- 0x06E4
		"00101100",	-- 0x06E5
		"00100000",	-- 0x06E6
		"01001100",	-- 0x06E7
		"00101000",	-- 0x06E8
		"01101111",	-- 0x06E9
		"01100001",	-- 0x06EA
		"01100100",	-- 0x06EB
		"00101001",	-- 0x06EC
		"00101100",	-- 0x06ED
		"00100000",	-- 0x06EE
		"01010010",	-- 0x06EF
		"00101000",	-- 0x06F0
		"01100101",	-- 0x06F1
		"01100111",	-- 0x06F2
		"01101001",	-- 0x06F3
		"01110011",	-- 0x06F4
		"01110100",	-- 0x06F5
		"01100101",	-- 0x06F6
		"01110010",	-- 0x06F7
		"00100000",	-- 0x06F8
		"01100100",	-- 0x06F9
		"01110101",	-- 0x06FA
		"01101101",	-- 0x06FB
		"01110000",	-- 0x06FC
		"00101001",	-- 0x06FD
		"00001101",	-- 0x06FE
		"00001010",	-- 0x06FF
		"00000000",	-- 0x0700
		"11110101",	-- 0x0701
		"11010101",	-- 0x0702
		"11100101",	-- 0x0703
		"00100001",	-- 0x0704
		"10000100",	-- 0x0705
		"00000111",	-- 0x0706
		"11001101",	-- 0x0707
		"01101001",	-- 0x0708
		"00001011",	-- 0x0709
		"11001101",	-- 0x070A
		"11100001",	-- 0x070B
		"00001010",	-- 0x070C
		"11111110",	-- 0x070D
		"00001101",	-- 0x070E
		"00101000",	-- 0x070F
		"11111001",	-- 0x0710
		"11111110",	-- 0x0711
		"00001010",	-- 0x0712
		"00101000",	-- 0x0713
		"11110101",	-- 0x0714
		"11111110",	-- 0x0715
		"00100000",	-- 0x0716
		"00101000",	-- 0x0717
		"11110001",	-- 0x0718
		"11001101",	-- 0x0719
		"10111001",	-- 0x071A
		"00001010",	-- 0x071B
		"11001101",	-- 0x071C
		"01100011",	-- 0x071D
		"00001011",	-- 0x071E
		"11111110",	-- 0x071F
		"00111010",	-- 0x0720
		"00100000",	-- 0x0721
		"01001110",	-- 0x0722
		"11001101",	-- 0x0723
		"11100111",	-- 0x0724
		"00001010",	-- 0x0725
		"01010111",	-- 0x0726
		"00011110",	-- 0x0727
		"00000000",	-- 0x0728
		"11001101",	-- 0x0729
		"01111110",	-- 0x072A
		"00000111",	-- 0x072B
		"11001101",	-- 0x072C
		"00001100",	-- 0x072D
		"00001011",	-- 0x072E
		"01111100",	-- 0x072F
		"11001101",	-- 0x0730
		"01111110",	-- 0x0731
		"00000111",	-- 0x0732
		"01111101",	-- 0x0733
		"11001101",	-- 0x0734
		"01111110",	-- 0x0735
		"00000111",	-- 0x0736
		"11001101",	-- 0x0737
		"11100111",	-- 0x0738
		"00001010",	-- 0x0739
		"11001101",	-- 0x073A
		"01111110",	-- 0x073B
		"00000111",	-- 0x073C
		"11111110",	-- 0x073D
		"00000001",	-- 0x073E
		"00100000",	-- 0x073F
		"00010010",	-- 0x0740
		"11001101",	-- 0x0741
		"11100111",	-- 0x0742
		"00001010",	-- 0x0743
		"11001101",	-- 0x0744
		"01111110",	-- 0x0745
		"00000111",	-- 0x0746
		"01111011",	-- 0x0747
		"10100111",	-- 0x0748
		"00101000",	-- 0x0749
		"00101100",	-- 0x074A
		"00100001",	-- 0x074B
		"10100100",	-- 0x074C
		"00000111",	-- 0x074D
		"11001101",	-- 0x074E
		"01101001",	-- 0x074F
		"00001011",	-- 0x0750
		"00011000",	-- 0x0751
		"00100100",	-- 0x0752
		"01111010",	-- 0x0753
		"10100111",	-- 0x0754
		"00101000",	-- 0x0755
		"00001011",	-- 0x0756
		"11001101",	-- 0x0757
		"11100111",	-- 0x0758
		"00001010",	-- 0x0759
		"11001101",	-- 0x075A
		"01111110",	-- 0x075B
		"00000111",	-- 0x075C
		"01110111",	-- 0x075D
		"00100011",	-- 0x075E
		"00010101",	-- 0x075F
		"00011000",	-- 0x0760
		"11110001",	-- 0x0761
		"11001101",	-- 0x0762
		"11100111",	-- 0x0763
		"00001010",	-- 0x0764
		"11001101",	-- 0x0765
		"01111110",	-- 0x0766
		"00000111",	-- 0x0767
		"01111011",	-- 0x0768
		"10100111",	-- 0x0769
		"00100000",	-- 0x076A
		"11011111",	-- 0x076B
		"11001101",	-- 0x076C
		"11010100",	-- 0x076D
		"00001010",	-- 0x076E
		"00011000",	-- 0x076F
		"10011001",	-- 0x0770
		"00100001",	-- 0x0771
		"10010101",	-- 0x0772
		"00000111",	-- 0x0773
		"11001101",	-- 0x0774
		"01101001",	-- 0x0775
		"00001011",	-- 0x0776
		"11001101",	-- 0x0777
		"11010100",	-- 0x0778
		"00001010",	-- 0x0779
		"11100001",	-- 0x077A
		"11010001",	-- 0x077B
		"11110001",	-- 0x077C
		"11001001",	-- 0x077D
		"01001111",	-- 0x077E
		"01111011",	-- 0x077F
		"10010001",	-- 0x0780
		"01011111",	-- 0x0781
		"01111001",	-- 0x0782
		"11001001",	-- 0x0783
		"01001001",	-- 0x0784
		"01001110",	-- 0x0785
		"01010100",	-- 0x0786
		"01000101",	-- 0x0787
		"01001100",	-- 0x0788
		"00100000",	-- 0x0789
		"01001000",	-- 0x078A
		"01000101",	-- 0x078B
		"01011000",	-- 0x078C
		"00100000",	-- 0x078D
		"01001100",	-- 0x078E
		"01001111",	-- 0x078F
		"01000001",	-- 0x0790
		"01000100",	-- 0x0791
		"00111010",	-- 0x0792
		"00100000",	-- 0x0793
		"00000000",	-- 0x0794
		"00100000",	-- 0x0795
		"01010011",	-- 0x0796
		"01111001",	-- 0x0797
		"01101110",	-- 0x0798
		"01110100",	-- 0x0799
		"01100001",	-- 0x079A
		"01111000",	-- 0x079B
		"00100000",	-- 0x079C
		"01100101",	-- 0x079D
		"01110010",	-- 0x079E
		"01110010",	-- 0x079F
		"01101111",	-- 0x07A0
		"01110010",	-- 0x07A1
		"00100001",	-- 0x07A2
		"00000000",	-- 0x07A3
		"00100000",	-- 0x07A4
		"01000011",	-- 0x07A5
		"01101000",	-- 0x07A6
		"01100101",	-- 0x07A7
		"01100011",	-- 0x07A8
		"01101011",	-- 0x07A9
		"01110011",	-- 0x07AA
		"01110101",	-- 0x07AB
		"01101101",	-- 0x07AC
		"00100000",	-- 0x07AD
		"01100101",	-- 0x07AE
		"01110010",	-- 0x07AF
		"01110010",	-- 0x07B0
		"01101111",	-- 0x07B1
		"01110010",	-- 0x07B2
		"00100001",	-- 0x07B3
		"00000000",	-- 0x07B4
		"11100101",	-- 0x07B5
		"00100001",	-- 0x07B6
		"11000100",	-- 0x07B7
		"00000111",	-- 0x07B8
		"11001101",	-- 0x07B9
		"01101001",	-- 0x07BA
		"00001011",	-- 0x07BB
		"00100001",	-- 0x07BC
		"01010011",	-- 0x07BD
		"00000001",	-- 0x07BE
		"11001101",	-- 0x07BF
		"01101001",	-- 0x07C0
		"00001011",	-- 0x07C1
		"11100001",	-- 0x07C2
		"11001001",	-- 0x07C3
		"01001001",	-- 0x07C4
		"01001110",	-- 0x07C5
		"01000110",	-- 0x07C6
		"01001111",	-- 0x07C7
		"00111010",	-- 0x07C8
		"00100000",	-- 0x07C9
		"00000000",	-- 0x07CA
		"11110101",	-- 0x07CB
		"11000101",	-- 0x07CC
		"11010101",	-- 0x07CD
		"11100101",	-- 0x07CE
		"00100001",	-- 0x07CF
		"00110110",	-- 0x07D0
		"00001000",	-- 0x07D1
		"11001101",	-- 0x07D2
		"01101001",	-- 0x07D3
		"00001011",	-- 0x07D4
		"11001101",	-- 0x07D5
		"00001100",	-- 0x07D6
		"00001011",	-- 0x07D7
		"11100101",	-- 0x07D8
		"10100111",	-- 0x07D9
		"00000001",	-- 0x07DA
		"00000000",	-- 0x07DB
		"10000000",	-- 0x07DC
		"11101101",	-- 0x07DD
		"01000010",	-- 0x07DE
		"11100001",	-- 0x07DF
		"00010001",	-- 0x07E0
		"00000000",	-- 0x07E1
		"00000000",	-- 0x07E2
		"00110000",	-- 0x07E3
		"00001000",	-- 0x07E4
		"00100001",	-- 0x07E5
		"01100111",	-- 0x07E6
		"00001000",	-- 0x07E7
		"11001101",	-- 0x07E8
		"01101001",	-- 0x07E9
		"00001011",	-- 0x07EA
		"00011000",	-- 0x07EB
		"00110110",	-- 0x07EC
		"00111110",	-- 0x07ED
		"00100000",	-- 0x07EE
		"11001101",	-- 0x07EF
		"01100011",	-- 0x07F0
		"00001011",	-- 0x07F1
		"11001101",	-- 0x07F2
		"11100001",	-- 0x07F3
		"00001010",	-- 0x07F4
		"11001101",	-- 0x07F5
		"10111001",	-- 0x07F6
		"00001010",	-- 0x07F7
		"11001101",	-- 0x07F8
		"10010001",	-- 0x07F9
		"00001010",	-- 0x07FA
		"00110000",	-- 0x07FB
		"00100110",	-- 0x07FC
		"11001101",	-- 0x07FD
		"10101110",	-- 0x07FE
		"00001010",	-- 0x07FF
		"11001101",	-- 0x0800
		"01000110",	-- 0x0801
		"00001011",	-- 0x0802
		"11001011",	-- 0x0803
		"00000111",	-- 0x0804
		"11001011",	-- 0x0805
		"00000111",	-- 0x0806
		"11001011",	-- 0x0807
		"00000111",	-- 0x0808
		"11001011",	-- 0x0809
		"00000111",	-- 0x080A
		"01000111",	-- 0x080B
		"11001101",	-- 0x080C
		"11100001",	-- 0x080D
		"00001010",	-- 0x080E
		"11001101",	-- 0x080F
		"10111001",	-- 0x0810
		"00001010",	-- 0x0811
		"11001101",	-- 0x0812
		"10010001",	-- 0x0813
		"00001010",	-- 0x0814
		"00110000",	-- 0x0815
		"00001100",	-- 0x0816
		"11001101",	-- 0x0817
		"10101110",	-- 0x0818
		"00001010",	-- 0x0819
		"11001101",	-- 0x081A
		"01000110",	-- 0x081B
		"00001011",	-- 0x081C
		"10110000",	-- 0x081D
		"01110111",	-- 0x081E
		"00100011",	-- 0x081F
		"00010011",	-- 0x0820
		"00011000",	-- 0x0821
		"11001010",	-- 0x0822
		"11001101",	-- 0x0823
		"11010100",	-- 0x0824
		"00001010",	-- 0x0825
		"01100010",	-- 0x0826
		"01101011",	-- 0x0827
		"11001101",	-- 0x0828
		"01010110",	-- 0x0829
		"00001011",	-- 0x082A
		"00100001",	-- 0x082B
		"01010110",	-- 0x082C
		"00001000",	-- 0x082D
		"11001101",	-- 0x082E
		"01101001",	-- 0x082F
		"00001011",	-- 0x0830
		"11100001",	-- 0x0831
		"11010001",	-- 0x0832
		"11000001",	-- 0x0833
		"11110001",	-- 0x0834
		"11001001",	-- 0x0835
		"01001100",	-- 0x0836
		"01001111",	-- 0x0837
		"01000001",	-- 0x0838
		"01000100",	-- 0x0839
		"00100000",	-- 0x083A
		"00101000",	-- 0x083B
		"01111000",	-- 0x083C
		"01111000",	-- 0x083D
		"00100000",	-- 0x083E
		"01101111",	-- 0x083F
		"01110010",	-- 0x0840
		"00100000",	-- 0x0841
		"01100101",	-- 0x0842
		"01101100",	-- 0x0843
		"01110011",	-- 0x0844
		"01100101",	-- 0x0845
		"00100000",	-- 0x0846
		"01110100",	-- 0x0847
		"01101111",	-- 0x0848
		"00100000",	-- 0x0849
		"01100101",	-- 0x084A
		"01101110",	-- 0x084B
		"01100100",	-- 0x084C
		"00101001",	-- 0x084D
		"00111010",	-- 0x084E
		"00100000",	-- 0x084F
		"01000001",	-- 0x0850
		"01000100",	-- 0x0851
		"01000100",	-- 0x0852
		"01010010",	-- 0x0853
		"00111101",	-- 0x0854
		"00000000",	-- 0x0855
		"00100000",	-- 0x0856
		"01100010",	-- 0x0857
		"01111001",	-- 0x0858
		"01110100",	-- 0x0859
		"01100101",	-- 0x085A
		"01110011",	-- 0x085B
		"00100000",	-- 0x085C
		"01101100",	-- 0x085D
		"01101111",	-- 0x085E
		"01100001",	-- 0x085F
		"01100100",	-- 0x0860
		"01100101",	-- 0x0861
		"01100100",	-- 0x0862
		"00101110",	-- 0x0863
		"00001101",	-- 0x0864
		"00001010",	-- 0x0865
		"00000000",	-- 0x0866
		"00100000",	-- 0x0867
		"01001001",	-- 0x0868
		"01101100",	-- 0x0869
		"01101100",	-- 0x086A
		"01100101",	-- 0x086B
		"01100111",	-- 0x086C
		"01100001",	-- 0x086D
		"01101100",	-- 0x086E
		"00100000",	-- 0x086F
		"01100001",	-- 0x0870
		"01100100",	-- 0x0871
		"01100100",	-- 0x0872
		"01110010",	-- 0x0873
		"01100101",	-- 0x0874
		"01110011",	-- 0x0875
		"01110011",	-- 0x0876
		"00100001",	-- 0x0877
		"00000000",	-- 0x0878
		"11110101",	-- 0x0879
		"11000101",	-- 0x087A
		"11010101",	-- 0x087B
		"11100101",	-- 0x087C
		"11111101",	-- 0x087D
		"11100101",	-- 0x087E
		"00100001",	-- 0x087F
		"11011000",	-- 0x0880
		"00001000",	-- 0x0881
		"11001101",	-- 0x0882
		"01101001",	-- 0x0883
		"00001011",	-- 0x0884
		"11001101",	-- 0x0885
		"00001100",	-- 0x0886
		"00001011",	-- 0x0887
		"00100010",	-- 0x0888
		"01011111",	-- 0x0889
		"11111011",	-- 0x088A
		"10100111",	-- 0x088B
		"00000001",	-- 0x088C
		"00000000",	-- 0x088D
		"10000000",	-- 0x088E
		"11101101",	-- 0x088F
		"01000010",	-- 0x0890
		"00110000",	-- 0x0891
		"00001000",	-- 0x0892
		"00100001",	-- 0x0893
		"11101001",	-- 0x0894
		"00001000",	-- 0x0895
		"11001101",	-- 0x0896
		"01101001",	-- 0x0897
		"00001011",	-- 0x0898
		"00011000",	-- 0x0899
		"00101000",	-- 0x089A
		"00100001",	-- 0x089B
		"00001100",	-- 0x089C
		"00001001",	-- 0x089D
		"11001101",	-- 0x089E
		"01101001",	-- 0x089F
		"00001011",	-- 0x08A0
		"00100001",	-- 0x08A1
		"01101101",	-- 0x08A2
		"11111011",	-- 0x08A3
		"00000110",	-- 0x08A4
		"01010001",	-- 0x08A5
		"11001101",	-- 0x08A6
		"00010111",	-- 0x08A7
		"00001011",	-- 0x08A8
		"11111101",	-- 0x08A9
		"00100001",	-- 0x08AA
		"10111110",	-- 0x08AB
		"11111011",	-- 0x08AC
		"00010001",	-- 0x08AD
		"01100001",	-- 0x08AE
		"11111011",	-- 0x08AF
		"11001101",	-- 0x08B0
		"00110101",	-- 0x08B1
		"00010000",	-- 0x08B2
		"00101010",	-- 0x08B3
		"01011111",	-- 0x08B4
		"11111011",	-- 0x08B5
		"00010001",	-- 0x08B6
		"00000000",	-- 0x08B7
		"00000000",	-- 0x08B8
		"11001101",	-- 0x08B9
		"01111010",	-- 0x08BA
		"00001101",	-- 0x08BB
		"00111000",	-- 0x08BC
		"00000101",	-- 0x08BD
		"01110111",	-- 0x08BE
		"00100011",	-- 0x08BF
		"00010011",	-- 0x08C0
		"00011000",	-- 0x08C1
		"11110110",	-- 0x08C2
		"11001101",	-- 0x08C3
		"11010100",	-- 0x08C4
		"00001010",	-- 0x08C5
		"01100010",	-- 0x08C6
		"01101011",	-- 0x08C7
		"11001101",	-- 0x08C8
		"01010110",	-- 0x08C9
		"00001011",	-- 0x08CA
		"00100001",	-- 0x08CB
		"11111011",	-- 0x08CC
		"00001000",	-- 0x08CD
		"11001101",	-- 0x08CE
		"01101001",	-- 0x08CF
		"00001011",	-- 0x08D0
		"11111101",	-- 0x08D1
		"11100001",	-- 0x08D2
		"11100001",	-- 0x08D3
		"11010001",	-- 0x08D4
		"11000001",	-- 0x08D5
		"11110001",	-- 0x08D6
		"11001001",	-- 0x08D7
		"01001100",	-- 0x08D8
		"01001111",	-- 0x08D9
		"01000001",	-- 0x08DA
		"01000100",	-- 0x08DB
		"00100000",	-- 0x08DC
		"01000110",	-- 0x08DD
		"01001001",	-- 0x08DE
		"01001100",	-- 0x08DF
		"01000101",	-- 0x08E0
		"00111010",	-- 0x08E1
		"00100000",	-- 0x08E2
		"01000001",	-- 0x08E3
		"01000100",	-- 0x08E4
		"01000100",	-- 0x08E5
		"01010010",	-- 0x08E6
		"00111101",	-- 0x08E7
		"00000000",	-- 0x08E8
		"00100000",	-- 0x08E9
		"01001001",	-- 0x08EA
		"01101100",	-- 0x08EB
		"01101100",	-- 0x08EC
		"01100101",	-- 0x08ED
		"01100111",	-- 0x08EE
		"01100001",	-- 0x08EF
		"01101100",	-- 0x08F0
		"00100000",	-- 0x08F1
		"01100001",	-- 0x08F2
		"01100100",	-- 0x08F3
		"01100100",	-- 0x08F4
		"01110010",	-- 0x08F5
		"01100101",	-- 0x08F6
		"01110011",	-- 0x08F7
		"01110011",	-- 0x08F8
		"00100001",	-- 0x08F9
		"00000000",	-- 0x08FA
		"00100000",	-- 0x08FB
		"01100010",	-- 0x08FC
		"01111001",	-- 0x08FD
		"01110100",	-- 0x08FE
		"01100101",	-- 0x08FF
		"01110011",	-- 0x0900
		"00100000",	-- 0x0901
		"01101100",	-- 0x0902
		"01101111",	-- 0x0903
		"01100001",	-- 0x0904
		"01100100",	-- 0x0905
		"01100101",	-- 0x0906
		"01100100",	-- 0x0907
		"00101110",	-- 0x0908
		"00001101",	-- 0x0909
		"00001010",	-- 0x090A
		"00000000",	-- 0x090B
		"00100000",	-- 0x090C
		"01000110",	-- 0x090D
		"01001001",	-- 0x090E
		"01001100",	-- 0x090F
		"01000101",	-- 0x0910
		"01001110",	-- 0x0911
		"01000001",	-- 0x0912
		"01001101",	-- 0x0913
		"01000101",	-- 0x0914
		"00111101",	-- 0x0915
		"00000000",	-- 0x0916
		"11100101",	-- 0x0917
		"00100001",	-- 0x0918
		"00100011",	-- 0x0919
		"00001001",	-- 0x091A
		"11001101",	-- 0x091B
		"01101001",	-- 0x091C
		"00001011",	-- 0x091D
		"11001101",	-- 0x091E
		"01100001",	-- 0x091F
		"00010011",	-- 0x0920
		"11100001",	-- 0x0921
		"11001001",	-- 0x0922
		"01001101",	-- 0x0923
		"01001111",	-- 0x0924
		"01010101",	-- 0x0925
		"01001110",	-- 0x0926
		"01010100",	-- 0x0927
		"00001101",	-- 0x0928
		"00001010",	-- 0x0929
		"00001101",	-- 0x092A
		"00001010",	-- 0x092B
		"00000000",	-- 0x092C
		"11110101",	-- 0x092D
		"11000101",	-- 0x092E
		"11010101",	-- 0x092F
		"11100101",	-- 0x0930
		"00100001",	-- 0x0931
		"01101101",	-- 0x0932
		"00001001",	-- 0x0933
		"11001101",	-- 0x0934
		"01101001",	-- 0x0935
		"00001011",	-- 0x0936
		"11001101",	-- 0x0937
		"00001100",	-- 0x0938
		"00001011",	-- 0x0939
		"11100101",	-- 0x093A
		"00100001",	-- 0x093B
		"01111001",	-- 0x093C
		"00001001",	-- 0x093D
		"11001101",	-- 0x093E
		"01101001",	-- 0x093F
		"00001011",	-- 0x0940
		"11001101",	-- 0x0941
		"00001100",	-- 0x0942
		"00001011",	-- 0x0943
		"01010100",	-- 0x0944
		"01011101",	-- 0x0945
		"10100111",	-- 0x0946
		"00000001",	-- 0x0947
		"00000000",	-- 0x0948
		"10000000",	-- 0x0949
		"11101101",	-- 0x094A
		"01000010",	-- 0x094B
		"00110000",	-- 0x094C
		"00001001",	-- 0x094D
		"00100001",	-- 0x094E
		"10000111",	-- 0x094F
		"00001001",	-- 0x0950
		"11001101",	-- 0x0951
		"01101001",	-- 0x0952
		"00001011",	-- 0x0953
		"11100001",	-- 0x0954
		"00011000",	-- 0x0955
		"00001110",	-- 0x0956
		"00100001",	-- 0x0957
		"01111110",	-- 0x0958
		"00001001",	-- 0x0959
		"11001101",	-- 0x095A
		"01101001",	-- 0x095B
		"00001011",	-- 0x095C
		"11001101",	-- 0x095D
		"00001100",	-- 0x095E
		"00001011",	-- 0x095F
		"01000100",	-- 0x0960
		"01001101",	-- 0x0961
		"11100001",	-- 0x0962
		"11101101",	-- 0x0963
		"10110000",	-- 0x0964
		"11001101",	-- 0x0965
		"11010100",	-- 0x0966
		"00001010",	-- 0x0967
		"11100001",	-- 0x0968
		"11010001",	-- 0x0969
		"11000001",	-- 0x096A
		"11110001",	-- 0x096B
		"11001001",	-- 0x096C
		"01001101",	-- 0x096D
		"01001111",	-- 0x096E
		"01010110",	-- 0x096F
		"01000101",	-- 0x0970
		"00111010",	-- 0x0971
		"00100000",	-- 0x0972
		"01000110",	-- 0x0973
		"01010010",	-- 0x0974
		"01001111",	-- 0x0975
		"01001101",	-- 0x0976
		"00111101",	-- 0x0977
		"00000000",	-- 0x0978
		"00100000",	-- 0x0979
		"01010100",	-- 0x097A
		"01001111",	-- 0x097B
		"00111101",	-- 0x097C
		"00000000",	-- 0x097D
		"00100000",	-- 0x097E
		"01001100",	-- 0x097F
		"01000101",	-- 0x0980
		"01001110",	-- 0x0981
		"01000111",	-- 0x0982
		"01010100",	-- 0x0983
		"01001000",	-- 0x0984
		"00111101",	-- 0x0985
		"00000000",	-- 0x0986
		"00100000",	-- 0x0987
		"01001001",	-- 0x0988
		"01101100",	-- 0x0989
		"01101100",	-- 0x098A
		"01100101",	-- 0x098B
		"01100111",	-- 0x098C
		"01100001",	-- 0x098D
		"01101100",	-- 0x098E
		"00100000",	-- 0x098F
		"01100100",	-- 0x0990
		"01100101",	-- 0x0991
		"01110011",	-- 0x0992
		"01110100",	-- 0x0993
		"01101001",	-- 0x0994
		"01101110",	-- 0x0995
		"01100001",	-- 0x0996
		"01110100",	-- 0x0997
		"01101001",	-- 0x0998
		"01101111",	-- 0x0999
		"01101110",	-- 0x099A
		"00100000",	-- 0x099B
		"01100001",	-- 0x099C
		"01100100",	-- 0x099D
		"01100100",	-- 0x099E
		"01110010",	-- 0x099F
		"01100101",	-- 0x09A0
		"01110011",	-- 0x09A1
		"01110011",	-- 0x09A2
		"00100001",	-- 0x09A3
		"00000000",	-- 0x09A4
		"11110101",	-- 0x09A5
		"11100101",	-- 0x09A6
		"00100001",	-- 0x09A7
		"11101100",	-- 0x09A8
		"00001001",	-- 0x09A9
		"11001101",	-- 0x09AA
		"01101001",	-- 0x09AB
		"00001011",	-- 0x09AC
		"11100001",	-- 0x09AD
		"11001101",	-- 0x09AE
		"00011101",	-- 0x09AF
		"00001010",	-- 0x09B0
		"11011001",	-- 0x09B1
		"00001000",	-- 0x09B2
		"11100101",	-- 0x09B3
		"00100001",	-- 0x09B4
		"00000011",	-- 0x09B5
		"00001010",	-- 0x09B6
		"11001101",	-- 0x09B7
		"01101001",	-- 0x09B8
		"00001011",	-- 0x09B9
		"11100001",	-- 0x09BA
		"11001101",	-- 0x09BB
		"00011101",	-- 0x09BC
		"00001010",	-- 0x09BD
		"00001000",	-- 0x09BE
		"11011001",	-- 0x09BF
		"11100101",	-- 0x09C0
		"00100001",	-- 0x09C1
		"00001001",	-- 0x09C2
		"00001010",	-- 0x09C3
		"11001101",	-- 0x09C4
		"01101001",	-- 0x09C5
		"00001011",	-- 0x09C6
		"11011101",	-- 0x09C7
		"11100101",	-- 0x09C8
		"11100001",	-- 0x09C9
		"11001101",	-- 0x09CA
		"01010110",	-- 0x09CB
		"00001011",	-- 0x09CC
		"00100001",	-- 0x09CD
		"00010011",	-- 0x09CE
		"00001010",	-- 0x09CF
		"11001101",	-- 0x09D0
		"01101001",	-- 0x09D1
		"00001011",	-- 0x09D2
		"11111101",	-- 0x09D3
		"11100101",	-- 0x09D4
		"11100001",	-- 0x09D5
		"11001101",	-- 0x09D6
		"01010110",	-- 0x09D7
		"00001011",	-- 0x09D8
		"00100001",	-- 0x09D9
		"00011000",	-- 0x09DA
		"00001010",	-- 0x09DB
		"11001101",	-- 0x09DC
		"01101001",	-- 0x09DD
		"00001011",	-- 0x09DE
		"00100001",	-- 0x09DF
		"00000000",	-- 0x09E0
		"00000000",	-- 0x09E1
		"00111001",	-- 0x09E2
		"11001101",	-- 0x09E3
		"01010110",	-- 0x09E4
		"00001011",	-- 0x09E5
		"11001101",	-- 0x09E6
		"11010100",	-- 0x09E7
		"00001010",	-- 0x09E8
		"11100001",	-- 0x09E9
		"11110001",	-- 0x09EA
		"11001001",	-- 0x09EB
		"01010010",	-- 0x09EC
		"01000101",	-- 0x09ED
		"01000111",	-- 0x09EE
		"01001001",	-- 0x09EF
		"01010011",	-- 0x09F0
		"01010100",	-- 0x09F1
		"01000101",	-- 0x09F2
		"01010010",	-- 0x09F3
		"00100000",	-- 0x09F4
		"01000100",	-- 0x09F5
		"01010101",	-- 0x09F6
		"01001101",	-- 0x09F7
		"01010000",	-- 0x09F8
		"00001101",	-- 0x09F9
		"00001010",	-- 0x09FA
		"00001101",	-- 0x09FB
		"00001010",	-- 0x09FC
		"00001001",	-- 0x09FD
		"00110001",	-- 0x09FE
		"01110011",	-- 0x09FF
		"01110100",	-- 0x0A00
		"00111010",	-- 0x0A01
		"00000000",	-- 0x0A02
		"00001001",	-- 0x0A03
		"00110010",	-- 0x0A04
		"01101110",	-- 0x0A05
		"01100100",	-- 0x0A06
		"00111010",	-- 0x0A07
		"00000000",	-- 0x0A08
		"00001001",	-- 0x0A09
		"01010000",	-- 0x0A0A
		"01010100",	-- 0x0A0B
		"01010010",	-- 0x0A0C
		"00111010",	-- 0x0A0D
		"00100000",	-- 0x0A0E
		"01001001",	-- 0x0A0F
		"01011000",	-- 0x0A10
		"00111101",	-- 0x0A11
		"00000000",	-- 0x0A12
		"00100000",	-- 0x0A13
		"01001001",	-- 0x0A14
		"01011001",	-- 0x0A15
		"00111101",	-- 0x0A16
		"00000000",	-- 0x0A17
		"00100000",	-- 0x0A18
		"01010011",	-- 0x0A19
		"01010000",	-- 0x0A1A
		"00111101",	-- 0x0A1B
		"00000000",	-- 0x0A1C
		"11100101",	-- 0x0A1D
		"00100001",	-- 0x0A1E
		"01001101",	-- 0x0A1F
		"00001010",	-- 0x0A20
		"11001101",	-- 0x0A21
		"01101001",	-- 0x0A22
		"00001011",	-- 0x0A23
		"11110101",	-- 0x0A24
		"11100001",	-- 0x0A25
		"11001101",	-- 0x0A26
		"01010110",	-- 0x0A27
		"00001011",	-- 0x0A28
		"00100001",	-- 0x0A29
		"01010010",	-- 0x0A2A
		"00001010",	-- 0x0A2B
		"11001101",	-- 0x0A2C
		"01101001",	-- 0x0A2D
		"00001011",	-- 0x0A2E
		"01100000",	-- 0x0A2F
		"01101001",	-- 0x0A30
		"11001101",	-- 0x0A31
		"01010110",	-- 0x0A32
		"00001011",	-- 0x0A33
		"00100001",	-- 0x0A34
		"01010111",	-- 0x0A35
		"00001010",	-- 0x0A36
		"11001101",	-- 0x0A37
		"01101001",	-- 0x0A38
		"00001011",	-- 0x0A39
		"01100010",	-- 0x0A3A
		"01101011",	-- 0x0A3B
		"11001101",	-- 0x0A3C
		"01010110",	-- 0x0A3D
		"00001011",	-- 0x0A3E
		"00100001",	-- 0x0A3F
		"01011100",	-- 0x0A40
		"00001010",	-- 0x0A41
		"11001101",	-- 0x0A42
		"01101001",	-- 0x0A43
		"00001011",	-- 0x0A44
		"11100001",	-- 0x0A45
		"11001101",	-- 0x0A46
		"01010110",	-- 0x0A47
		"00001011",	-- 0x0A48
		"11001101",	-- 0x0A49
		"11010100",	-- 0x0A4A
		"00001010",	-- 0x0A4B
		"11001001",	-- 0x0A4C
		"00100000",	-- 0x0A4D
		"01000001",	-- 0x0A4E
		"01000110",	-- 0x0A4F
		"00111101",	-- 0x0A50
		"00000000",	-- 0x0A51
		"00100000",	-- 0x0A52
		"01000010",	-- 0x0A53
		"01000011",	-- 0x0A54
		"00111101",	-- 0x0A55
		"00000000",	-- 0x0A56
		"00100000",	-- 0x0A57
		"01000100",	-- 0x0A58
		"01000101",	-- 0x0A59
		"00111101",	-- 0x0A5A
		"00000000",	-- 0x0A5B
		"00100000",	-- 0x0A5C
		"01001000",	-- 0x0A5D
		"01001100",	-- 0x0A5E
		"00111101",	-- 0x0A5F
		"00000000",	-- 0x0A60
		"00100001",	-- 0x0A61
		"01101110",	-- 0x0A62
		"00001010",	-- 0x0A63
		"11001101",	-- 0x0A64
		"01101001",	-- 0x0A65
		"00001011",	-- 0x0A66
		"11001101",	-- 0x0A67
		"00001100",	-- 0x0A68
		"00001011",	-- 0x0A69
		"11001101",	-- 0x0A6A
		"11010100",	-- 0x0A6B
		"00001010",	-- 0x0A6C
		"11101001",	-- 0x0A6D
		"01010011",	-- 0x0A6E
		"01010100",	-- 0x0A6F
		"01000001",	-- 0x0A70
		"01010010",	-- 0x0A71
		"01010100",	-- 0x0A72
		"00111010",	-- 0x0A73
		"00100000",	-- 0x0A74
		"01000001",	-- 0x0A75
		"01000100",	-- 0x0A76
		"01000100",	-- 0x0A77
		"01010010",	-- 0x0A78
		"00111101",	-- 0x0A79
		"00000000",	-- 0x0A7A
		"11100101",	-- 0x0A7B
		"00100001",	-- 0x0A7C
		"10000111",	-- 0x0A7D
		"00001010",	-- 0x0A7E
		"11001101",	-- 0x0A7F
		"01101001",	-- 0x0A80
		"00001011",	-- 0x0A81
		"11001101",	-- 0x0A82
		"01011001",	-- 0x0A83
		"00010110",	-- 0x0A84
		"11100001",	-- 0x0A85
		"11001001",	-- 0x0A86
		"01010101",	-- 0x0A87
		"01001110",	-- 0x0A88
		"01001101",	-- 0x0A89
		"01001111",	-- 0x0A8A
		"01010101",	-- 0x0A8B
		"01001110",	-- 0x0A8C
		"01010100",	-- 0x0A8D
		"00001101",	-- 0x0A8E
		"00001010",	-- 0x0A8F
		"00000000",	-- 0x0A90
		"11111110",	-- 0x0A91
		"01000111",	-- 0x0A92
		"11010000",	-- 0x0A93
		"11111110",	-- 0x0A94
		"00110000",	-- 0x0A95
		"00110000",	-- 0x0A96
		"00000010",	-- 0x0A97
		"00111111",	-- 0x0A98
		"11001001",	-- 0x0A99
		"11111110",	-- 0x0A9A
		"00111010",	-- 0x0A9B
		"11011000",	-- 0x0A9C
		"11111110",	-- 0x0A9D
		"01000001",	-- 0x0A9E
		"00110000",	-- 0x0A9F
		"00000010",	-- 0x0AA0
		"00111111",	-- 0x0AA1
		"11001001",	-- 0x0AA2
		"00110111",	-- 0x0AA3
		"11001001",	-- 0x0AA4
		"11111110",	-- 0x0AA5
		"00100000",	-- 0x0AA6
		"00110000",	-- 0x0AA7
		"00000010",	-- 0x0AA8
		"00111111",	-- 0x0AA9
		"11001001",	-- 0x0AAA
		"11111110",	-- 0x0AAB
		"01111111",	-- 0x0AAC
		"11001001",	-- 0x0AAD
		"11111110",	-- 0x0AAE
		"00111010",	-- 0x0AAF
		"00111000",	-- 0x0AB0
		"00000010",	-- 0x0AB1
		"11010110",	-- 0x0AB2
		"00000111",	-- 0x0AB3
		"11010110",	-- 0x0AB4
		"00110000",	-- 0x0AB5
		"11100110",	-- 0x0AB6
		"00001111",	-- 0x0AB7
		"11001001",	-- 0x0AB8
		"11111110",	-- 0x0AB9
		"01100001",	-- 0x0ABA
		"11011000",	-- 0x0ABB
		"11111110",	-- 0x0ABC
		"01111011",	-- 0x0ABD
		"11010000",	-- 0x0ABE
		"11100110",	-- 0x0ABF
		"01011111",	-- 0x0AC0
		"11001001",	-- 0x0AC1
		"11010101",	-- 0x0AC2
		"11100101",	-- 0x0AC3
		"00011010",	-- 0x0AC4
		"11111110",	-- 0x0AC5
		"00000000",	-- 0x0AC6
		"00101000",	-- 0x0AC7
		"00000111",	-- 0x0AC8
		"10111110",	-- 0x0AC9
		"00100000",	-- 0x0ACA
		"00000100",	-- 0x0ACB
		"00100011",	-- 0x0ACC
		"00010011",	-- 0x0ACD
		"00011000",	-- 0x0ACE
		"11110100",	-- 0x0ACF
		"10010110",	-- 0x0AD0
		"11100001",	-- 0x0AD1
		"11010001",	-- 0x0AD2
		"11001001",	-- 0x0AD3
		"11110101",	-- 0x0AD4
		"00111110",	-- 0x0AD5
		"00001101",	-- 0x0AD6
		"11001101",	-- 0x0AD7
		"01100011",	-- 0x0AD8
		"00001011",	-- 0x0AD9
		"00111110",	-- 0x0ADA
		"00001010",	-- 0x0ADB
		"11001101",	-- 0x0ADC
		"01100011",	-- 0x0ADD
		"00001011",	-- 0x0ADE
		"11110001",	-- 0x0ADF
		"11001001",	-- 0x0AE0
		"11001101",	-- 0x0AE1
		"01111001",	-- 0x0AE2
		"00001011",	-- 0x0AE3
		"11011011",	-- 0x0AE4
		"00000000",	-- 0x0AE5
		"11001001",	-- 0x0AE6
		"11000101",	-- 0x0AE7
		"11001101",	-- 0x0AE8
		"11111010",	-- 0x0AE9
		"00001010",	-- 0x0AEA
		"11001011",	-- 0x0AEB
		"00000111",	-- 0x0AEC
		"11001011",	-- 0x0AED
		"00000111",	-- 0x0AEE
		"11001011",	-- 0x0AEF
		"00000111",	-- 0x0AF0
		"11001011",	-- 0x0AF1
		"00000111",	-- 0x0AF2
		"01000111",	-- 0x0AF3
		"11001101",	-- 0x0AF4
		"11111010",	-- 0x0AF5
		"00001010",	-- 0x0AF6
		"10110000",	-- 0x0AF7
		"11000001",	-- 0x0AF8
		"11001001",	-- 0x0AF9
		"11001101",	-- 0x0AFA
		"11100001",	-- 0x0AFB
		"00001010",	-- 0x0AFC
		"11001101",	-- 0x0AFD
		"10111001",	-- 0x0AFE
		"00001010",	-- 0x0AFF
		"11001101",	-- 0x0B00
		"10010001",	-- 0x0B01
		"00001010",	-- 0x0B02
		"00110000",	-- 0x0B03
		"11110101",	-- 0x0B04
		"11001101",	-- 0x0B05
		"10101110",	-- 0x0B06
		"00001010",	-- 0x0B07
		"11001101",	-- 0x0B08
		"01000110",	-- 0x0B09
		"00001011",	-- 0x0B0A
		"11001001",	-- 0x0B0B
		"11110101",	-- 0x0B0C
		"11001101",	-- 0x0B0D
		"11100111",	-- 0x0B0E
		"00001010",	-- 0x0B0F
		"01100111",	-- 0x0B10
		"11001101",	-- 0x0B11
		"11100111",	-- 0x0B12
		"00001010",	-- 0x0B13
		"01101111",	-- 0x0B14
		"11110001",	-- 0x0B15
		"11001001",	-- 0x0B16
		"11110101",	-- 0x0B17
		"11000101",	-- 0x0B18
		"11100101",	-- 0x0B19
		"11001101",	-- 0x0B1A
		"11100001",	-- 0x0B1B
		"00001010",	-- 0x0B1C
		"11111110",	-- 0x0B1D
		"00001101",	-- 0x0B1E
		"00101000",	-- 0x0B1F
		"11111001",	-- 0x0B20
		"11001101",	-- 0x0B21
		"10111001",	-- 0x0B22
		"00001010",	-- 0x0B23
		"11001101",	-- 0x0B24
		"01100011",	-- 0x0B25
		"00001011",	-- 0x0B26
		"11111110",	-- 0x0B27
		"00001010",	-- 0x0B28
		"00101000",	-- 0x0B29
		"00000100",	-- 0x0B2A
		"01110111",	-- 0x0B2B
		"00100011",	-- 0x0B2C
		"00010000",	-- 0x0B2D
		"11101011",	-- 0x0B2E
		"00110110",	-- 0x0B2F
		"00000000",	-- 0x0B30
		"11100001",	-- 0x0B31
		"11000001",	-- 0x0B32
		"11110001",	-- 0x0B33
		"11001001",	-- 0x0B34
		"11110101",	-- 0x0B35
		"11000101",	-- 0x0B36
		"01000111",	-- 0x0B37
		"00001111",	-- 0x0B38
		"00001111",	-- 0x0B39
		"00001111",	-- 0x0B3A
		"00001111",	-- 0x0B3B
		"11001101",	-- 0x0B3C
		"01000110",	-- 0x0B3D
		"00001011",	-- 0x0B3E
		"01111000",	-- 0x0B3F
		"11001101",	-- 0x0B40
		"01000110",	-- 0x0B41
		"00001011",	-- 0x0B42
		"11000001",	-- 0x0B43
		"11110001",	-- 0x0B44
		"11001001",	-- 0x0B45
		"11110101",	-- 0x0B46
		"11100110",	-- 0x0B47
		"00001111",	-- 0x0B48
		"11000110",	-- 0x0B49
		"00110000",	-- 0x0B4A
		"11111110",	-- 0x0B4B
		"00111010",	-- 0x0B4C
		"00111000",	-- 0x0B4D
		"00000010",	-- 0x0B4E
		"11000110",	-- 0x0B4F
		"00000111",	-- 0x0B50
		"11001101",	-- 0x0B51
		"01100011",	-- 0x0B52
		"00001011",	-- 0x0B53
		"11110001",	-- 0x0B54
		"11001001",	-- 0x0B55
		"11100101",	-- 0x0B56
		"11110101",	-- 0x0B57
		"01111100",	-- 0x0B58
		"11001101",	-- 0x0B59
		"00110101",	-- 0x0B5A
		"00001011",	-- 0x0B5B
		"01111101",	-- 0x0B5C
		"11001101",	-- 0x0B5D
		"00110101",	-- 0x0B5E
		"00001011",	-- 0x0B5F
		"11110001",	-- 0x0B60
		"11100001",	-- 0x0B61
		"11001001",	-- 0x0B62
		"11001101",	-- 0x0B63
		"10000010",	-- 0x0B64
		"00001011",	-- 0x0B65
		"11010011",	-- 0x0B66
		"00000000",	-- 0x0B67
		"11001001",	-- 0x0B68
		"11110101",	-- 0x0B69
		"11100101",	-- 0x0B6A
		"01111110",	-- 0x0B6B
		"11111110",	-- 0x0B6C
		"00000000",	-- 0x0B6D
		"00101000",	-- 0x0B6E
		"00000110",	-- 0x0B6F
		"11001101",	-- 0x0B70
		"01100011",	-- 0x0B71
		"00001011",	-- 0x0B72
		"00100011",	-- 0x0B73
		"00011000",	-- 0x0B74
		"11110101",	-- 0x0B75
		"11100001",	-- 0x0B76
		"11110001",	-- 0x0B77
		"11001001",	-- 0x0B78
		"11110101",	-- 0x0B79
		"11011011",	-- 0x0B7A
		"00000101",	-- 0x0B7B
		"11001011",	-- 0x0B7C
		"01000111",	-- 0x0B7D
		"00101000",	-- 0x0B7E
		"11111010",	-- 0x0B7F
		"11110001",	-- 0x0B80
		"11001001",	-- 0x0B81
		"11110101",	-- 0x0B82
		"11011011",	-- 0x0B83
		"00000101",	-- 0x0B84
		"11001011",	-- 0x0B85
		"01101111",	-- 0x0B86
		"00101000",	-- 0x0B87
		"11111010",	-- 0x0B88
		"11110001",	-- 0x0B89
		"11001001",	-- 0x0B8A
		"11110101",	-- 0x0B8B
		"11000101",	-- 0x0B8C
		"11100101",	-- 0x0B8D
		"11001101",	-- 0x0B8E
		"11110001",	-- 0x0B8F
		"00001100",	-- 0x0B90
		"00111000",	-- 0x0B91
		"00101110",	-- 0x0B92
		"00111110",	-- 0x0B93
		"10100000",	-- 0x0B94
		"11010011",	-- 0x0B95
		"00010111",	-- 0x0B96
		"11001101",	-- 0x0B97
		"11110001",	-- 0x0B98
		"00001100",	-- 0x0B99
		"00111000",	-- 0x0B9A
		"00100101",	-- 0x0B9B
		"00111110",	-- 0x0B9C
		"11101100",	-- 0x0B9D
		"11010011",	-- 0x0B9E
		"00010111",	-- 0x0B9F
		"11001101",	-- 0x0BA0
		"11110001",	-- 0x0BA1
		"00001100",	-- 0x0BA2
		"00111000",	-- 0x0BA3
		"00011100",	-- 0x0BA4
		"11001101",	-- 0x0BA5
		"00100010",	-- 0x0BA6
		"00001100",	-- 0x0BA7
		"00111000",	-- 0x0BA8
		"00010111",	-- 0x0BA9
		"11001101",	-- 0x0BAA
		"11100001",	-- 0x0BAB
		"00001011",	-- 0x0BAC
		"00111000",	-- 0x0BAD
		"00010010",	-- 0x0BAE
		"00100001",	-- 0x0BAF
		"00000000",	-- 0x0BB0
		"11111110",	-- 0x0BB1
		"00000110",	-- 0x0BB2
		"00000000",	-- 0x0BB3
		"11011011",	-- 0x0BB4
		"00010000",	-- 0x0BB5
		"01001111",	-- 0x0BB6
		"11011011",	-- 0x0BB7
		"00011000",	-- 0x0BB8
		"01110111",	-- 0x0BB9
		"00100011",	-- 0x0BBA
		"01110001",	-- 0x0BBB
		"00100011",	-- 0x0BBC
		"00010000",	-- 0x0BBD
		"11110101",	-- 0x0BBE
		"00011000",	-- 0x0BBF
		"00000110",	-- 0x0BC0
		"00100001",	-- 0x0BC1
		"11001011",	-- 0x0BC2
		"00001011",	-- 0x0BC3
		"11001101",	-- 0x0BC4
		"01101001",	-- 0x0BC5
		"00001011",	-- 0x0BC6
		"11100001",	-- 0x0BC7
		"11000001",	-- 0x0BC8
		"11110001",	-- 0x0BC9
		"11001001",	-- 0x0BCA
		"01000110",	-- 0x0BCB
		"01000001",	-- 0x0BCC
		"01010100",	-- 0x0BCD
		"01000001",	-- 0x0BCE
		"01001100",	-- 0x0BCF
		"00101000",	-- 0x0BD0
		"01001001",	-- 0x0BD1
		"01000100",	-- 0x0BD2
		"01000101",	-- 0x0BD3
		"00101001",	-- 0x0BD4
		"00111010",	-- 0x0BD5
		"00100000",	-- 0x0BD6
		"01000001",	-- 0x0BD7
		"01100010",	-- 0x0BD8
		"01101111",	-- 0x0BD9
		"01110010",	-- 0x0BDA
		"01110100",	-- 0x0BDB
		"01100101",	-- 0x0BDC
		"01100100",	-- 0x0BDD
		"00100001",	-- 0x0BDE
		"00001101",	-- 0x0BDF
		"00001010",	-- 0x0BE0
		"11000101",	-- 0x0BE1
		"10100111",	-- 0x0BE2
		"00000110",	-- 0x0BE3
		"11111111",	-- 0x0BE4
		"11011011",	-- 0x0BE5
		"00010111",	-- 0x0BE6
		"11001011",	-- 0x0BE7
		"01011111",	-- 0x0BE8
		"00100000",	-- 0x0BE9
		"00010000",	-- 0x0BEA
		"11000101",	-- 0x0BEB
		"00000110",	-- 0x0BEC
		"00000000",	-- 0x0BED
		"00000000",	-- 0x0BEE
		"00010000",	-- 0x0BEF
		"11111101",	-- 0x0BF0
		"11000001",	-- 0x0BF1
		"00010000",	-- 0x0BF2
		"11110001",	-- 0x0BF3
		"00110111",	-- 0x0BF4
		"00100001",	-- 0x0BF5
		"11111101",	-- 0x0BF6
		"00001011",	-- 0x0BF7
		"11001101",	-- 0x0BF8
		"01101001",	-- 0x0BF9
		"00001011",	-- 0x0BFA
		"11000001",	-- 0x0BFB
		"11001001",	-- 0x0BFC
		"01000110",	-- 0x0BFD
		"01000001",	-- 0x0BFE
		"01010100",	-- 0x0BFF
		"01000001",	-- 0x0C00
		"01001100",	-- 0x0C01
		"00101000",	-- 0x0C02
		"01001001",	-- 0x0C03
		"01000100",	-- 0x0C04
		"01000101",	-- 0x0C05
		"00101001",	-- 0x0C06
		"00111010",	-- 0x0C07
		"00100000",	-- 0x0C08
		"01101001",	-- 0x0C09
		"01100100",	-- 0x0C0A
		"01100101",	-- 0x0C0B
		"01011111",	-- 0x0C0C
		"01100010",	-- 0x0C0D
		"01100110",	-- 0x0C0E
		"01110010",	-- 0x0C0F
		"01011111",	-- 0x0C10
		"01110010",	-- 0x0C11
		"01100101",	-- 0x0C12
		"01100001",	-- 0x0C13
		"01100100",	-- 0x0C14
		"01111001",	-- 0x0C15
		"00100000",	-- 0x0C16
		"01110100",	-- 0x0C17
		"01101001",	-- 0x0C18
		"01101101",	-- 0x0C19
		"01100101",	-- 0x0C1A
		"01101111",	-- 0x0C1B
		"01110101",	-- 0x0C1C
		"01110100",	-- 0x0C1D
		"00100001",	-- 0x0C1E
		"00001101",	-- 0x0C1F
		"00001010",	-- 0x0C20
		"00000000",	-- 0x0C21
		"10100111",	-- 0x0C22
		"11011011",	-- 0x0C23
		"00010111",	-- 0x0C24
		"11001011",	-- 0x0C25
		"01000111",	-- 0x0C26
		"00101000",	-- 0x0C27
		"00000001",	-- 0x0C28
		"00110111",	-- 0x0C29
		"11001001",	-- 0x0C2A
		"11000101",	-- 0x0C2B
		"11100101",	-- 0x0C2C
		"11001101",	-- 0x0C2D
		"11110001",	-- 0x0C2E
		"00001100",	-- 0x0C2F
		"00111000",	-- 0x0C30
		"00101001",	-- 0x0C31
		"11001101",	-- 0x0C32
		"11011010",	-- 0x0C33
		"00001100",	-- 0x0C34
		"11001101",	-- 0x0C35
		"11110001",	-- 0x0C36
		"00001100",	-- 0x0C37
		"00111000",	-- 0x0C38
		"00100001",	-- 0x0C39
		"00111110",	-- 0x0C3A
		"00100000",	-- 0x0C3B
		"11010011",	-- 0x0C3C
		"00010111",	-- 0x0C3D
		"11001101",	-- 0x0C3E
		"11110001",	-- 0x0C3F
		"00001100",	-- 0x0C40
		"00111000",	-- 0x0C41
		"00011000",	-- 0x0C42
		"11001101",	-- 0x0C43
		"00100010",	-- 0x0C44
		"00001100",	-- 0x0C45
		"00111000",	-- 0x0C46
		"00010011",	-- 0x0C47
		"11001101",	-- 0x0C48
		"11100001",	-- 0x0C49
		"00001011",	-- 0x0C4A
		"00111000",	-- 0x0C4B
		"00001110",	-- 0x0C4C
		"00000110",	-- 0x0C4D
		"00000000",	-- 0x0C4E
		"11011011",	-- 0x0C4F
		"00010000",	-- 0x0C50
		"01110111",	-- 0x0C51
		"00100011",	-- 0x0C52
		"11011011",	-- 0x0C53
		"00011000",	-- 0x0C54
		"01110111",	-- 0x0C55
		"00100011",	-- 0x0C56
		"00010000",	-- 0x0C57
		"11110110",	-- 0x0C58
		"00011000",	-- 0x0C59
		"00000110",	-- 0x0C5A
		"00100001",	-- 0x0C5B
		"01100100",	-- 0x0C5C
		"00001100",	-- 0x0C5D
		"11001101",	-- 0x0C5E
		"01101001",	-- 0x0C5F
		"00001011",	-- 0x0C60
		"11100001",	-- 0x0C61
		"11000001",	-- 0x0C62
		"11001001",	-- 0x0C63
		"01000110",	-- 0x0C64
		"01000001",	-- 0x0C65
		"01010100",	-- 0x0C66
		"01000001",	-- 0x0C67
		"01001100",	-- 0x0C68
		"00101000",	-- 0x0C69
		"01001001",	-- 0x0C6A
		"01000100",	-- 0x0C6B
		"01000101",	-- 0x0C6C
		"00101001",	-- 0x0C6D
		"00111010",	-- 0x0C6E
		"00100000",	-- 0x0C6F
		"01101001",	-- 0x0C70
		"01100100",	-- 0x0C71
		"01100101",	-- 0x0C72
		"01011111",	-- 0x0C73
		"01110010",	-- 0x0C74
		"01110011",	-- 0x0C75
		"00100000",	-- 0x0C76
		"01110100",	-- 0x0C77
		"01101001",	-- 0x0C78
		"01101101",	-- 0x0C79
		"01100101",	-- 0x0C7A
		"01101111",	-- 0x0C7B
		"01110101",	-- 0x0C7C
		"01110100",	-- 0x0C7D
		"00100001",	-- 0x0C7E
		"00001101",	-- 0x0C7F
		"00001010",	-- 0x0C80
		"00000000",	-- 0x0C81
		"11000101",	-- 0x0C82
		"11100101",	-- 0x0C83
		"11001101",	-- 0x0C84
		"11110001",	-- 0x0C85
		"00001100",	-- 0x0C86
		"00111000",	-- 0x0C87
		"00101010",	-- 0x0C88
		"11001101",	-- 0x0C89
		"11011010",	-- 0x0C8A
		"00001100",	-- 0x0C8B
		"11001101",	-- 0x0C8C
		"11110001",	-- 0x0C8D
		"00001100",	-- 0x0C8E
		"00111000",	-- 0x0C8F
		"00100010",	-- 0x0C90
		"00111110",	-- 0x0C91
		"00110000",	-- 0x0C92
		"11010011",	-- 0x0C93
		"00010111",	-- 0x0C94
		"11001101",	-- 0x0C95
		"11110001",	-- 0x0C96
		"00001100",	-- 0x0C97
		"00111000",	-- 0x0C98
		"00011001",	-- 0x0C99
		"11001101",	-- 0x0C9A
		"00100010",	-- 0x0C9B
		"00001100",	-- 0x0C9C
		"00111000",	-- 0x0C9D
		"00010100",	-- 0x0C9E
		"11001101",	-- 0x0C9F
		"11100001",	-- 0x0CA0
		"00001011",	-- 0x0CA1
		"00111000",	-- 0x0CA2
		"00001111",	-- 0x0CA3
		"00000110",	-- 0x0CA4
		"00000000",	-- 0x0CA5
		"01111110",	-- 0x0CA6
		"01001111",	-- 0x0CA7
		"00100011",	-- 0x0CA8
		"01111110",	-- 0x0CA9
		"11010011",	-- 0x0CAA
		"00011000",	-- 0x0CAB
		"01111001",	-- 0x0CAC
		"11010011",	-- 0x0CAD
		"00010000",	-- 0x0CAE
		"00010000",	-- 0x0CAF
		"11110101",	-- 0x0CB0
		"00011000",	-- 0x0CB1
		"00000110",	-- 0x0CB2
		"00100001",	-- 0x0CB3
		"10111100",	-- 0x0CB4
		"00001100",	-- 0x0CB5
		"11001101",	-- 0x0CB6
		"01101001",	-- 0x0CB7
		"00001011",	-- 0x0CB8
		"11100001",	-- 0x0CB9
		"11000001",	-- 0x0CBA
		"11001001",	-- 0x0CBB
		"01000110",	-- 0x0CBC
		"01000001",	-- 0x0CBD
		"01010100",	-- 0x0CBE
		"01000001",	-- 0x0CBF
		"01001100",	-- 0x0CC0
		"00101000",	-- 0x0CC1
		"01001001",	-- 0x0CC2
		"01000100",	-- 0x0CC3
		"01000101",	-- 0x0CC4
		"00101001",	-- 0x0CC5
		"00111010",	-- 0x0CC6
		"00100000",	-- 0x0CC7
		"01101001",	-- 0x0CC8
		"01100100",	-- 0x0CC9
		"01100101",	-- 0x0CCA
		"01011111",	-- 0x0CCB
		"01110111",	-- 0x0CCC
		"01110011",	-- 0x0CCD
		"00100000",	-- 0x0CCE
		"01110100",	-- 0x0CCF
		"01101001",	-- 0x0CD0
		"01101101",	-- 0x0CD1
		"01100101",	-- 0x0CD2
		"01101111",	-- 0x0CD3
		"01110101",	-- 0x0CD4
		"01110100",	-- 0x0CD5
		"00100001",	-- 0x0CD6
		"00001101",	-- 0x0CD7
		"00001010",	-- 0x0CD8
		"00000000",	-- 0x0CD9
		"11110101",	-- 0x0CDA
		"00111110",	-- 0x0CDB
		"00000001",	-- 0x0CDC
		"11010011",	-- 0x0CDD
		"00010010",	-- 0x0CDE
		"01111011",	-- 0x0CDF
		"11010011",	-- 0x0CE0
		"00010011",	-- 0x0CE1
		"01111010",	-- 0x0CE2
		"11010011",	-- 0x0CE3
		"00010100",	-- 0x0CE4
		"01111001",	-- 0x0CE5
		"11010011",	-- 0x0CE6
		"00010101",	-- 0x0CE7
		"01111000",	-- 0x0CE8
		"11100110",	-- 0x0CE9
		"00001111",	-- 0x0CEA
		"11110110",	-- 0x0CEB
		"11100000",	-- 0x0CEC
		"11010011",	-- 0x0CED
		"00010110",	-- 0x0CEE
		"11110001",	-- 0x0CEF
		"11001001",	-- 0x0CF0
		"11000101",	-- 0x0CF1
		"10100111",	-- 0x0CF2
		"00000110",	-- 0x0CF3
		"11111111",	-- 0x0CF4
		"11011011",	-- 0x0CF5
		"00010111",	-- 0x0CF6
		"11100110",	-- 0x0CF7
		"11000000",	-- 0x0CF8
		"11101110",	-- 0x0CF9
		"01000000",	-- 0x0CFA
		"00101000",	-- 0x0CFB
		"00010101",	-- 0x0CFC
		"11000101",	-- 0x0CFD
		"00000110",	-- 0x0CFE
		"00000000",	-- 0x0CFF
		"00000000",	-- 0x0D00
		"00010000",	-- 0x0D01
		"11111101",	-- 0x0D02
		"11000001",	-- 0x0D03
		"00010000",	-- 0x0D04
		"11101111",	-- 0x0D05
		"00110111",	-- 0x0D06
		"00100001",	-- 0x0D07
		"00010100",	-- 0x0D08
		"00001101",	-- 0x0D09
		"11001101",	-- 0x0D0A
		"01101001",	-- 0x0D0B
		"00001011",	-- 0x0D0C
		"11011011",	-- 0x0D0D
		"00010001",	-- 0x0D0E
		"11001101",	-- 0x0D0F
		"00110101",	-- 0x0D10
		"00001011",	-- 0x0D11
		"11000001",	-- 0x0D12
		"11001001",	-- 0x0D13
		"01000110",	-- 0x0D14
		"01000001",	-- 0x0D15
		"01010100",	-- 0x0D16
		"01000001",	-- 0x0D17
		"01001100",	-- 0x0D18
		"00101000",	-- 0x0D19
		"01001001",	-- 0x0D1A
		"01000100",	-- 0x0D1B
		"01000101",	-- 0x0D1C
		"00101001",	-- 0x0D1D
		"00111010",	-- 0x0D1E
		"00100000",	-- 0x0D1F
		"01101001",	-- 0x0D20
		"01100100",	-- 0x0D21
		"01100101",	-- 0x0D22
		"01011111",	-- 0x0D23
		"01110010",	-- 0x0D24
		"01100101",	-- 0x0D25
		"01100001",	-- 0x0D26
		"01100100",	-- 0x0D27
		"01111001",	-- 0x0D28
		"00100000",	-- 0x0D29
		"01110100",	-- 0x0D2A
		"01101001",	-- 0x0D2B
		"01101101",	-- 0x0D2C
		"01100101",	-- 0x0D2D
		"01101111",	-- 0x0D2E
		"01110101",	-- 0x0D2F
		"01110100",	-- 0x0D30
		"00100001",	-- 0x0D31
		"00001101",	-- 0x0D32
		"00001010",	-- 0x0D33
		"00000000",	-- 0x0D34
		"00100001",	-- 0x0D35
		"01001100",	-- 0x0D36
		"11111011",	-- 0x0D37
		"00110110",	-- 0x0D38
		"00000000",	-- 0x0D39
		"00100001",	-- 0x0D3A
		"01000110",	-- 0x0D3B
		"00001101",	-- 0x0D3C
		"11001101",	-- 0x0D3D
		"01101001",	-- 0x0D3E
		"00001011",	-- 0x0D3F
		"00111110",	-- 0x0D40
		"00000000",	-- 0x0D41
		"00110010",	-- 0x0D42
		"11111111",	-- 0x0D43
		"11111111",	-- 0x0D44
		"11000111",	-- 0x0D45
		"01000011",	-- 0x0D46
		"01001100",	-- 0x0D47
		"01000101",	-- 0x0D48
		"01000001",	-- 0x0D49
		"01010010",	-- 0x0D4A
		"00001101",	-- 0x0D4B
		"00001010",	-- 0x0D4C
		"00000000",	-- 0x0D4D
		"00011001",	-- 0x0D4E
		"11011001",	-- 0x0D4F
		"11101101",	-- 0x0D50
		"01011010",	-- 0x0D51
		"11011001",	-- 0x0D52
		"11001001",	-- 0x0D53
		"10100111",	-- 0x0D54
		"11101101",	-- 0x0D55
		"01100010",	-- 0x0D56
		"11011001",	-- 0x0D57
		"11101101",	-- 0x0D58
		"01100010",	-- 0x0D59
		"01111000",	-- 0x0D5A
		"00000110",	-- 0x0D5B
		"00100000",	-- 0x0D5C
		"11001011",	-- 0x0D5D
		"00101111",	-- 0x0D5E
		"11001011",	-- 0x0D5F
		"00011001",	-- 0x0D60
		"11011001",	-- 0x0D61
		"11001011",	-- 0x0D62
		"00011000",	-- 0x0D63
		"11001011",	-- 0x0D64
		"00011001",	-- 0x0D65
		"00110000",	-- 0x0D66
		"00000101",	-- 0x0D67
		"00011001",	-- 0x0D68
		"11011001",	-- 0x0D69
		"11101101",	-- 0x0D6A
		"01011010",	-- 0x0D6B
		"11011001",	-- 0x0D6C
		"11001011",	-- 0x0D6D
		"00100011",	-- 0x0D6E
		"11001011",	-- 0x0D6F
		"00010010",	-- 0x0D70
		"11011001",	-- 0x0D71
		"11001011",	-- 0x0D72
		"00010011",	-- 0x0D73
		"11001011",	-- 0x0D74
		"00010010",	-- 0x0D75
		"00010000",	-- 0x0D76
		"11100101",	-- 0x0D77
		"11011001",	-- 0x0D78
		"11001001",	-- 0x0D79
		"11000101",	-- 0x0D7A
		"11010101",	-- 0x0D7B
		"11100101",	-- 0x0D7C
		"11111101",	-- 0x0D7D
		"01111110",	-- 0x0D7E
		"00001100",	-- 0x0D7F
		"11111101",	-- 0x0D80
		"10111110",	-- 0x0D81
		"00010011",	-- 0x0D82
		"00100000",	-- 0x0D83
		"00011100",	-- 0x0D84
		"11111101",	-- 0x0D85
		"01111110",	-- 0x0D86
		"00001101",	-- 0x0D87
		"11111101",	-- 0x0D88
		"10111110",	-- 0x0D89
		"00010100",	-- 0x0D8A
		"00100000",	-- 0x0D8B
		"00010100",	-- 0x0D8C
		"11111101",	-- 0x0D8D
		"01111110",	-- 0x0D8E
		"00001110",	-- 0x0D8F
		"11111101",	-- 0x0D90
		"10111110",	-- 0x0D91
		"00010101",	-- 0x0D92
		"00100000",	-- 0x0D93
		"00001100",	-- 0x0D94
		"11111101",	-- 0x0D95
		"01111110",	-- 0x0D96
		"00001111",	-- 0x0D97
		"11111101",	-- 0x0D98
		"10111110",	-- 0x0D99
		"00010110",	-- 0x0D9A
		"00100000",	-- 0x0D9B
		"00000100",	-- 0x0D9C
		"00110111",	-- 0x0D9D
		"11000011",	-- 0x0D9E
		"10001010",	-- 0x0D9F
		"00001110",	-- 0x0DA0
		"11111101",	-- 0x0DA1
		"01111110",	-- 0x0DA2
		"00010011",	-- 0x0DA3
		"11111110",	-- 0x0DA4
		"00000000",	-- 0x0DA5
		"11000010",	-- 0x0DA6
		"01010110",	-- 0x0DA7
		"00001110",	-- 0x0DA8
		"11111101",	-- 0x0DA9
		"01111110",	-- 0x0DAA
		"00010100",	-- 0x0DAB
		"11100110",	-- 0x0DAC
		"00000001",	-- 0x0DAD
		"11000010",	-- 0x0DAE
		"01010110",	-- 0x0DAF
		"00001110",	-- 0x0DB0
		"11111101",	-- 0x0DB1
		"01111110",	-- 0x0DB2
		"00010111",	-- 0x0DB3
		"11111110",	-- 0x0DB4
		"00000000",	-- 0x0DB5
		"00100000",	-- 0x0DB6
		"00010101",	-- 0x0DB7
		"11111101",	-- 0x0DB8
		"01111110",	-- 0x0DB9
		"00011000",	-- 0x0DBA
		"11111110",	-- 0x0DBB
		"00000000",	-- 0x0DBC
		"00100000",	-- 0x0DBD
		"00001110",	-- 0x0DBE
		"11111101",	-- 0x0DBF
		"01111110",	-- 0x0DC0
		"00010000",	-- 0x0DC1
		"11111101",	-- 0x0DC2
		"01110111",	-- 0x0DC3
		"00010111",	-- 0x0DC4
		"11111101",	-- 0x0DC5
		"01111110",	-- 0x0DC6
		"00010001",	-- 0x0DC7
		"11111101",	-- 0x0DC8
		"01110111",	-- 0x0DC9
		"00011000",	-- 0x0DCA
		"00011000",	-- 0x0DCB
		"00110111",	-- 0x0DCC
		"11111101",	-- 0x0DCD
		"01111110",	-- 0x0DCE
		"00011101",	-- 0x0DCF
		"00100000",	-- 0x0DD0
		"01000011",	-- 0x0DD1
		"00101010",	-- 0x0DD2
		"11110100",	-- 0x0DD3
		"11111101",	-- 0x0DD4
		"11111101",	-- 0x0DD5
		"01001110",	-- 0x0DD6
		"00011000",	-- 0x0DD7
		"00000110",	-- 0x0DD8
		"00000000",	-- 0x0DD9
		"00001001",	-- 0x0DDA
		"01010100",	-- 0x0DDB
		"01011101",	-- 0x0DDC
		"00000001",	-- 0x0DDD
		"00000000",	-- 0x0DDE
		"00000000",	-- 0x0DDF
		"00101010",	-- 0x0DE0
		"11110110",	-- 0x0DE1
		"11111101",	-- 0x0DE2
		"11101101",	-- 0x0DE3
		"01001010",	-- 0x0DE4
		"01000100",	-- 0x0DE5
		"01001101",	-- 0x0DE6
		"00100001",	-- 0x0DE7
		"00000000",	-- 0x0DE8
		"11111110",	-- 0x0DE9
		"11001101",	-- 0x0DEA
		"00101011",	-- 0x0DEB
		"00001100",	-- 0x0DEC
		"00000110",	-- 0x0DED
		"00000000",	-- 0x0DEE
		"11111101",	-- 0x0DEF
		"01001110",	-- 0x0DF0
		"00010111",	-- 0x0DF1
		"11001011",	-- 0x0DF2
		"00100001",	-- 0x0DF3
		"11001011",	-- 0x0DF4
		"00010000",	-- 0x0DF5
		"00100001",	-- 0x0DF6
		"00000000",	-- 0x0DF7
		"11111110",	-- 0x0DF8
		"00001001",	-- 0x0DF9
		"01001110",	-- 0x0DFA
		"00100011",	-- 0x0DFB
		"01000110",	-- 0x0DFC
		"00101011",	-- 0x0DFD
		"11111101",	-- 0x0DFE
		"01110001",	-- 0x0DFF
		"00010111",	-- 0x0E00
		"11111101",	-- 0x0E01
		"01110000",	-- 0x0E02
		"00010111",	-- 0x0E03
		"00111010",	-- 0x0E04
		"11100101",	-- 0x0E05
		"11111101",	-- 0x0E06
		"11111101",	-- 0x0E07
		"01110111",	-- 0x0E08
		"00011101",	-- 0x0E09
		"11111101",	-- 0x0E0A
		"01101110",	-- 0x0E0B
		"00010111",	-- 0x0E0C
		"11111101",	-- 0x0E0D
		"01100110",	-- 0x0E0E
		"00011000",	-- 0x0E0F
		"11001101",	-- 0x0E10
		"01001111",	-- 0x0E11
		"00010001",	-- 0x0E12
		"00011000",	-- 0x0E13
		"00100110",	-- 0x0E14
		"10100111",	-- 0x0E15
		"00000001",	-- 0x0E16
		"00000001",	-- 0x0E17
		"00000000",	-- 0x0E18
		"11111101",	-- 0x0E19
		"01101110",	-- 0x0E1A
		"00011001",	-- 0x0E1B
		"11111101",	-- 0x0E1C
		"01100110",	-- 0x0E1D
		"00011010",	-- 0x0E1E
		"00001001",	-- 0x0E1F
		"11111101",	-- 0x0E20
		"01110101",	-- 0x0E21
		"00011001",	-- 0x0E22
		"01011101",	-- 0x0E23
		"11111101",	-- 0x0E24
		"01110100",	-- 0x0E25
		"00011010",	-- 0x0E26
		"01010100",	-- 0x0E27
		"11111101",	-- 0x0E28
		"01101110",	-- 0x0E29
		"00011011",	-- 0x0E2A
		"11111101",	-- 0x0E2B
		"01100110",	-- 0x0E2C
		"00011100",	-- 0x0E2D
		"00000001",	-- 0x0E2E
		"00000000",	-- 0x0E2F
		"00000000",	-- 0x0E30
		"11101101",	-- 0x0E31
		"01001010",	-- 0x0E32
		"11111101",	-- 0x0E33
		"01110101",	-- 0x0E34
		"00011011",	-- 0x0E35
		"01001101",	-- 0x0E36
		"11111101",	-- 0x0E37
		"01110100",	-- 0x0E38
		"00011100",	-- 0x0E39
		"01000100",	-- 0x0E3A
		"11111101",	-- 0x0E3B
		"01110011",	-- 0x0E3C
		"00011001",	-- 0x0E3D
		"11111101",	-- 0x0E3E
		"01110010",	-- 0x0E3F
		"00011010",	-- 0x0E40
		"11111101",	-- 0x0E41
		"01110001",	-- 0x0E42
		"00011011",	-- 0x0E43
		"11111101",	-- 0x0E44
		"01110000",	-- 0x0E45
		"00011100",	-- 0x0E46
		"11111101",	-- 0x0E47
		"11100101",	-- 0x0E48
		"11100001",	-- 0x0E49
		"11000101",	-- 0x0E4A
		"00000001",	-- 0x0E4B
		"00011110",	-- 0x0E4C
		"00000000",	-- 0x0E4D
		"00001001",	-- 0x0E4E
		"11000001",	-- 0x0E4F
		"11001101",	-- 0x0E50
		"00101011",	-- 0x0E51
		"00001100",	-- 0x0E52
		"11111101",	-- 0x0E53
		"00110101",	-- 0x0E54
		"00011101",	-- 0x0E55
		"11111101",	-- 0x0E56
		"11100101",	-- 0x0E57
		"11100001",	-- 0x0E58
		"00000001",	-- 0x0E59
		"00011110",	-- 0x0E5A
		"00000000",	-- 0x0E5B
		"00001001",	-- 0x0E5C
		"11111101",	-- 0x0E5D
		"01001110",	-- 0x0E5E
		"00010011",	-- 0x0E5F
		"11111101",	-- 0x0E60
		"01111110",	-- 0x0E61
		"00010100",	-- 0x0E62
		"11100110",	-- 0x0E63
		"00000001",	-- 0x0E64
		"01000111",	-- 0x0E65
		"00001001",	-- 0x0E66
		"01111110",	-- 0x0E67
		"11111101",	-- 0x0E68
		"01101110",	-- 0x0E69
		"00010011",	-- 0x0E6A
		"11111101",	-- 0x0E6B
		"01100110",	-- 0x0E6C
		"00010100",	-- 0x0E6D
		"00000001",	-- 0x0E6E
		"00000001",	-- 0x0E6F
		"00000000",	-- 0x0E70
		"00001001",	-- 0x0E71
		"11111101",	-- 0x0E72
		"01110101",	-- 0x0E73
		"00010011",	-- 0x0E74
		"11111101",	-- 0x0E75
		"01110100",	-- 0x0E76
		"00010100",	-- 0x0E77
		"00000001",	-- 0x0E78
		"00000000",	-- 0x0E79
		"00000000",	-- 0x0E7A
		"11111101",	-- 0x0E7B
		"01101110",	-- 0x0E7C
		"00010101",	-- 0x0E7D
		"11111101",	-- 0x0E7E
		"01100110",	-- 0x0E7F
		"00010110",	-- 0x0E80
		"11101101",	-- 0x0E81
		"01001010",	-- 0x0E82
		"11111101",	-- 0x0E83
		"01110101",	-- 0x0E84
		"00010101",	-- 0x0E85
		"11111101",	-- 0x0E86
		"01110100",	-- 0x0E87
		"00010110",	-- 0x0E88
		"10100111",	-- 0x0E89
		"11100001",	-- 0x0E8A
		"11010001",	-- 0x0E8B
		"11000001",	-- 0x0E8C
		"11001001",	-- 0x0E8D
		"11110101",	-- 0x0E8E
		"11000101",	-- 0x0E8F
		"11010101",	-- 0x0E90
		"11100101",	-- 0x0E91
		"00111110",	-- 0x0E92
		"00000000",	-- 0x0E93
		"11111101",	-- 0x0E94
		"11100101",	-- 0x0E95
		"11100001",	-- 0x0E96
		"01110111",	-- 0x0E97
		"01010100",	-- 0x0E98
		"01011101",	-- 0x0E99
		"00010011",	-- 0x0E9A
		"00000001",	-- 0x0E9B
		"00011110",	-- 0x0E9C
		"00000000",	-- 0x0E9D
		"11101101",	-- 0x0E9E
		"10110000",	-- 0x0E9F
		"11100001",	-- 0x0EA0
		"11010001",	-- 0x0EA1
		"11000001",	-- 0x0EA2
		"11110001",	-- 0x0EA3
		"11001001",	-- 0x0EA4
		"11110101",	-- 0x0EA5
		"11100101",	-- 0x0EA6
		"00100001",	-- 0x0EA7
		"00110111",	-- 0x0EA8
		"00001111",	-- 0x0EA9
		"11001101",	-- 0x0EAA
		"01101001",	-- 0x0EAB
		"00001011",	-- 0x0EAC
		"11111101",	-- 0x0EAD
		"11100101",	-- 0x0EAE
		"11100001",	-- 0x0EAF
		"11001101",	-- 0x0EB0
		"01010110",	-- 0x0EB1
		"00001011",	-- 0x0EB2
		"00100001",	-- 0x0EB3
		"01010000",	-- 0x0EB4
		"00001111",	-- 0x0EB5
		"11001101",	-- 0x0EB6
		"01101001",	-- 0x0EB7
		"00001011",	-- 0x0EB8
		"11111101",	-- 0x0EB9
		"11100101",	-- 0x0EBA
		"11100001",	-- 0x0EBB
		"11001101",	-- 0x0EBC
		"01101001",	-- 0x0EBD
		"00001011",	-- 0x0EBE
		"00100001",	-- 0x0EBF
		"01100101",	-- 0x0EC0
		"00001111",	-- 0x0EC1
		"11001101",	-- 0x0EC2
		"01101001",	-- 0x0EC3
		"00001011",	-- 0x0EC4
		"11111101",	-- 0x0EC5
		"01100110",	-- 0x0EC6
		"00001111",	-- 0x0EC7
		"11111101",	-- 0x0EC8
		"01101110",	-- 0x0EC9
		"00001110",	-- 0x0ECA
		"11001101",	-- 0x0ECB
		"01010110",	-- 0x0ECC
		"00001011",	-- 0x0ECD
		"11111101",	-- 0x0ECE
		"01100110",	-- 0x0ECF
		"00001101",	-- 0x0ED0
		"11111101",	-- 0x0ED1
		"01101110",	-- 0x0ED2
		"00001100",	-- 0x0ED3
		"11001101",	-- 0x0ED4
		"01010110",	-- 0x0ED5
		"00001011",	-- 0x0ED6
		"00100001",	-- 0x0ED7
		"01111010",	-- 0x0ED8
		"00001111",	-- 0x0ED9
		"11001101",	-- 0x0EDA
		"01101001",	-- 0x0EDB
		"00001011",	-- 0x0EDC
		"11111101",	-- 0x0EDD
		"01100110",	-- 0x0EDE
		"00010001",	-- 0x0EDF
		"11111101",	-- 0x0EE0
		"01101110",	-- 0x0EE1
		"00010000",	-- 0x0EE2
		"11001101",	-- 0x0EE3
		"01010110",	-- 0x0EE4
		"00001011",	-- 0x0EE5
		"00100001",	-- 0x0EE6
		"10001111",	-- 0x0EE7
		"00001111",	-- 0x0EE8
		"11001101",	-- 0x0EE9
		"01101001",	-- 0x0EEA
		"00001011",	-- 0x0EEB
		"11111101",	-- 0x0EEC
		"01111110",	-- 0x0EED
		"00010010",	-- 0x0EEE
		"11001101",	-- 0x0EEF
		"00110101",	-- 0x0EF0
		"00001011",	-- 0x0EF1
		"00100001",	-- 0x0EF2
		"10100100",	-- 0x0EF3
		"00001111",	-- 0x0EF4
		"11001101",	-- 0x0EF5
		"01101001",	-- 0x0EF6
		"00001011",	-- 0x0EF7
		"11111101",	-- 0x0EF8
		"01100110",	-- 0x0EF9
		"00010110",	-- 0x0EFA
		"11111101",	-- 0x0EFB
		"01101110",	-- 0x0EFC
		"00010101",	-- 0x0EFD
		"11001101",	-- 0x0EFE
		"01010110",	-- 0x0EFF
		"00001011",	-- 0x0F00
		"11111101",	-- 0x0F01
		"01100110",	-- 0x0F02
		"00010100",	-- 0x0F03
		"11111101",	-- 0x0F04
		"01101110",	-- 0x0F05
		"00010011",	-- 0x0F06
		"11001101",	-- 0x0F07
		"01010110",	-- 0x0F08
		"00001011",	-- 0x0F09
		"00100001",	-- 0x0F0A
		"10111001",	-- 0x0F0B
		"00001111",	-- 0x0F0C
		"11001101",	-- 0x0F0D
		"01101001",	-- 0x0F0E
		"00001011",	-- 0x0F0F
		"11111101",	-- 0x0F10
		"01100110",	-- 0x0F11
		"00011000",	-- 0x0F12
		"11111101",	-- 0x0F13
		"01101110",	-- 0x0F14
		"00010111",	-- 0x0F15
		"11001101",	-- 0x0F16
		"01010110",	-- 0x0F17
		"00001011",	-- 0x0F18
		"00100001",	-- 0x0F19
		"11001110",	-- 0x0F1A
		"00001111",	-- 0x0F1B
		"11001101",	-- 0x0F1C
		"01101001",	-- 0x0F1D
		"00001011",	-- 0x0F1E
		"11111101",	-- 0x0F1F
		"01100110",	-- 0x0F20
		"00011100",	-- 0x0F21
		"11111101",	-- 0x0F22
		"01101110",	-- 0x0F23
		"00011011",	-- 0x0F24
		"11001101",	-- 0x0F25
		"01010110",	-- 0x0F26
		"00001011",	-- 0x0F27
		"11111101",	-- 0x0F28
		"01100110",	-- 0x0F29
		"00011010",	-- 0x0F2A
		"11111101",	-- 0x0F2B
		"01101110",	-- 0x0F2C
		"00011001",	-- 0x0F2D
		"11001101",	-- 0x0F2E
		"01010110",	-- 0x0F2F
		"00001011",	-- 0x0F30
		"11001101",	-- 0x0F31
		"11010100",	-- 0x0F32
		"00001010",	-- 0x0F33
		"11100001",	-- 0x0F34
		"11110001",	-- 0x0F35
		"11001001",	-- 0x0F36
		"01000100",	-- 0x0F37
		"01110101",	-- 0x0F38
		"01101101",	-- 0x0F39
		"01110000",	-- 0x0F3A
		"00100000",	-- 0x0F3B
		"01101111",	-- 0x0F3C
		"01100110",	-- 0x0F3D
		"00100000",	-- 0x0F3E
		"01000110",	-- 0x0F3F
		"01000011",	-- 0x0F40
		"01000010",	-- 0x0F41
		"00100000",	-- 0x0F42
		"01100001",	-- 0x0F43
		"01110100",	-- 0x0F44
		"00100000",	-- 0x0F45
		"01100001",	-- 0x0F46
		"01100100",	-- 0x0F47
		"01100100",	-- 0x0F48
		"01110010",	-- 0x0F49
		"01100101",	-- 0x0F4A
		"01110011",	-- 0x0F4B
		"01110011",	-- 0x0F4C
		"00111010",	-- 0x0F4D
		"00100000",	-- 0x0F4E
		"00000000",	-- 0x0F4F
		"00001101",	-- 0x0F50
		"00001010",	-- 0x0F51
		"00001001",	-- 0x0F52
		"01000110",	-- 0x0F53
		"01101001",	-- 0x0F54
		"01101100",	-- 0x0F55
		"01100101",	-- 0x0F56
		"00100000",	-- 0x0F57
		"01101110",	-- 0x0F58
		"01100001",	-- 0x0F59
		"01101101",	-- 0x0F5A
		"01100101",	-- 0x0F5B
		"00100000",	-- 0x0F5C
		"00100000",	-- 0x0F5D
		"00100000",	-- 0x0F5E
		"00100000",	-- 0x0F5F
		"00100000",	-- 0x0F60
		"00100000",	-- 0x0F61
		"00111010",	-- 0x0F62
		"00100000",	-- 0x0F63
		"00000000",	-- 0x0F64
		"00001101",	-- 0x0F65
		"00001010",	-- 0x0F66
		"00001001",	-- 0x0F67
		"01000110",	-- 0x0F68
		"01101001",	-- 0x0F69
		"01101100",	-- 0x0F6A
		"01100101",	-- 0x0F6B
		"00100000",	-- 0x0F6C
		"01110011",	-- 0x0F6D
		"01101001",	-- 0x0F6E
		"01111010",	-- 0x0F6F
		"01100101",	-- 0x0F70
		"00100000",	-- 0x0F71
		"00100000",	-- 0x0F72
		"00100000",	-- 0x0F73
		"00100000",	-- 0x0F74
		"00100000",	-- 0x0F75
		"00100000",	-- 0x0F76
		"00111010",	-- 0x0F77
		"00100000",	-- 0x0F78
		"00000000",	-- 0x0F79
		"00001101",	-- 0x0F7A
		"00001010",	-- 0x0F7B
		"00001001",	-- 0x0F7C
		"00110001",	-- 0x0F7D
		"01110011",	-- 0x0F7E
		"01110100",	-- 0x0F7F
		"00100000",	-- 0x0F80
		"01100011",	-- 0x0F81
		"01101100",	-- 0x0F82
		"01110101",	-- 0x0F83
		"01110011",	-- 0x0F84
		"01110100",	-- 0x0F85
		"01100101",	-- 0x0F86
		"01110010",	-- 0x0F87
		"00100000",	-- 0x0F88
		"00100000",	-- 0x0F89
		"00100000",	-- 0x0F8A
		"00100000",	-- 0x0F8B
		"00111010",	-- 0x0F8C
		"00100000",	-- 0x0F8D
		"00000000",	-- 0x0F8E
		"00001101",	-- 0x0F8F
		"00001010",	-- 0x0F90
		"00001001",	-- 0x0F91
		"01000110",	-- 0x0F92
		"01101001",	-- 0x0F93
		"01101100",	-- 0x0F94
		"01100101",	-- 0x0F95
		"00100000",	-- 0x0F96
		"01110100",	-- 0x0F97
		"01111001",	-- 0x0F98
		"01110000",	-- 0x0F99
		"01100101",	-- 0x0F9A
		"00100000",	-- 0x0F9B
		"00100000",	-- 0x0F9C
		"00100000",	-- 0x0F9D
		"00100000",	-- 0x0F9E
		"00100000",	-- 0x0F9F
		"00100000",	-- 0x0FA0
		"00111010",	-- 0x0FA1
		"00100000",	-- 0x0FA2
		"00000000",	-- 0x0FA3
		"00001101",	-- 0x0FA4
		"00001010",	-- 0x0FA5
		"00001001",	-- 0x0FA6
		"01000110",	-- 0x0FA7
		"01101001",	-- 0x0FA8
		"01101100",	-- 0x0FA9
		"01100101",	-- 0x0FAA
		"00100000",	-- 0x0FAB
		"01110000",	-- 0x0FAC
		"01101111",	-- 0x0FAD
		"01101001",	-- 0x0FAE
		"01101110",	-- 0x0FAF
		"01110100",	-- 0x0FB0
		"01100101",	-- 0x0FB1
		"01110010",	-- 0x0FB2
		"00100000",	-- 0x0FB3
		"00100000",	-- 0x0FB4
		"00100000",	-- 0x0FB5
		"00111010",	-- 0x0FB6
		"00100000",	-- 0x0FB7
		"00000000",	-- 0x0FB8
		"00001101",	-- 0x0FB9
		"00001010",	-- 0x0FBA
		"00001001",	-- 0x0FBB
		"01000011",	-- 0x0FBC
		"01110101",	-- 0x0FBD
		"01110010",	-- 0x0FBE
		"01110010",	-- 0x0FBF
		"01100101",	-- 0x0FC0
		"01101110",	-- 0x0FC1
		"01110100",	-- 0x0FC2
		"00100000",	-- 0x0FC3
		"01100011",	-- 0x0FC4
		"01101100",	-- 0x0FC5
		"01110101",	-- 0x0FC6
		"01110011",	-- 0x0FC7
		"01110100",	-- 0x0FC8
		"01100101",	-- 0x0FC9
		"01110010",	-- 0x0FCA
		"00111010",	-- 0x0FCB
		"00100000",	-- 0x0FCC
		"00000000",	-- 0x0FCD
		"00001101",	-- 0x0FCE
		"00001010",	-- 0x0FCF
		"00001001",	-- 0x0FD0
		"01000011",	-- 0x0FD1
		"01110101",	-- 0x0FD2
		"01110010",	-- 0x0FD3
		"01110010",	-- 0x0FD4
		"01100101",	-- 0x0FD5
		"01101110",	-- 0x0FD6
		"01110100",	-- 0x0FD7
		"00100000",	-- 0x0FD8
		"01110011",	-- 0x0FD9
		"01100101",	-- 0x0FDA
		"01100011",	-- 0x0FDB
		"01110100",	-- 0x0FDC
		"01101111",	-- 0x0FDD
		"01110010",	-- 0x0FDE
		"00100000",	-- 0x0FDF
		"00111010",	-- 0x0FE0
		"00100000",	-- 0x0FE1
		"00000000",	-- 0x0FE2
		"11110101",	-- 0x0FE3
		"11000101",	-- 0x0FE4
		"11010101",	-- 0x0FE5
		"11100101",	-- 0x0FE6
		"11101101",	-- 0x0FE7
		"01010011",	-- 0x0FE8
		"01011101",	-- 0x0FE9
		"11111011",	-- 0x0FEA
		"00111110",	-- 0x0FEB
		"00100000",	-- 0x0FEC
		"00000110",	-- 0x0FED
		"00001011",	-- 0x0FEE
		"00010010",	-- 0x0FEF
		"00010011",	-- 0x0FF0
		"00010000",	-- 0x0FF1
		"11111100",	-- 0x0FF2
		"00111110",	-- 0x0FF3
		"00000000",	-- 0x0FF4
		"00010010",	-- 0x0FF5
		"11101101",	-- 0x0FF6
		"01011011",	-- 0x0FF7
		"01011101",	-- 0x0FF8
		"11111011",	-- 0x0FF9
		"00000110",	-- 0x0FFA
		"00001000",	-- 0x0FFB
		"01111110",	-- 0x0FFC
		"11111110",	-- 0x0FFD
		"00000000",	-- 0x0FFE
		"00101000",	-- 0x0FFF
		"00101111",	-- 0x1000
		"11111110",	-- 0x1001
		"00101110",	-- 0x1002
		"00101000",	-- 0x1003
		"00010010",	-- 0x1004
		"00010010",	-- 0x1005
		"00010011",	-- 0x1006
		"00100011",	-- 0x1007
		"00000101",	-- 0x1008
		"00100000",	-- 0x1009
		"11110001",	-- 0x100A
		"01111110",	-- 0x100B
		"11111110",	-- 0x100C
		"00000000",	-- 0x100D
		"00101000",	-- 0x100E
		"00100000",	-- 0x100F
		"11111110",	-- 0x1010
		"00101110",	-- 0x1011
		"00101000",	-- 0x1012
		"00000011",	-- 0x1013
		"00100011",	-- 0x1014
		"00011000",	-- 0x1015
		"11110100",	-- 0x1016
		"00100011",	-- 0x1017
		"11100101",	-- 0x1018
		"00101010",	-- 0x1019
		"01011101",	-- 0x101A
		"11111011",	-- 0x101B
		"00000001",	-- 0x101C
		"00001000",	-- 0x101D
		"00000000",	-- 0x101E
		"00001001",	-- 0x101F
		"01010100",	-- 0x1020
		"01011101",	-- 0x1021
		"11100001",	-- 0x1022
		"00000110",	-- 0x1023
		"00000011",	-- 0x1024
		"01111110",	-- 0x1025
		"11111110",	-- 0x1026
		"00000000",	-- 0x1027
		"00101000",	-- 0x1028
		"00000110",	-- 0x1029
		"00010010",	-- 0x102A
		"00010011",	-- 0x102B
		"00100011",	-- 0x102C
		"00000101",	-- 0x102D
		"00100000",	-- 0x102E
		"11110101",	-- 0x102F
		"11100001",	-- 0x1030
		"11010001",	-- 0x1031
		"11000001",	-- 0x1032
		"11110001",	-- 0x1033
		"11001001",	-- 0x1034
		"11110101",	-- 0x1035
		"11000101",	-- 0x1036
		"11010101",	-- 0x1037
		"11011101",	-- 0x1038
		"11100101",	-- 0x1039
		"00100010",	-- 0x103A
		"01010101",	-- 0x103B
		"11111011",	-- 0x103C
		"00100001",	-- 0x103D
		"11011100",	-- 0x103E
		"11111101",	-- 0x103F
		"01111110",	-- 0x1040
		"11111110",	-- 0x1041
		"00000000",	-- 0x1042
		"11001010",	-- 0x1043
		"11101100",	-- 0x1044
		"00010000",	-- 0x1045
		"11001101",	-- 0x1046
		"10001110",	-- 0x1047
		"00001110",	-- 0x1048
		"11111101",	-- 0x1049
		"11100101",	-- 0x104A
		"11010001",	-- 0x104B
		"00101010",	-- 0x104C
		"01010101",	-- 0x104D
		"11111011",	-- 0x104E
		"11001101",	-- 0x104F
		"11100011",	-- 0x1050
		"00001111",	-- 0x1051
		"00100001",	-- 0x1052
		"00000000",	-- 0x1053
		"11111110",	-- 0x1054
		"00000001",	-- 0x1055
		"00000000",	-- 0x1056
		"00000010",	-- 0x1057
		"00001001",	-- 0x1058
		"00100010",	-- 0x1059
		"01011011",	-- 0x105A
		"11111011",	-- 0x105B
		"00101010",	-- 0x105C
		"11111000",	-- 0x105D
		"11111101",	-- 0x105E
		"00100010",	-- 0x105F
		"01010111",	-- 0x1060
		"11111011",	-- 0x1061
		"00101010",	-- 0x1062
		"11111010",	-- 0x1063
		"11111101",	-- 0x1064
		"00100010",	-- 0x1065
		"01011001",	-- 0x1066
		"11111011",	-- 0x1067
		"11101101",	-- 0x1068
		"01001011",	-- 0x1069
		"01011001",	-- 0x106A
		"11111011",	-- 0x106B
		"11101101",	-- 0x106C
		"01011011",	-- 0x106D
		"01010111",	-- 0x106E
		"11111011",	-- 0x106F
		"00100001",	-- 0x1070
		"00000000",	-- 0x1071
		"11111110",	-- 0x1072
		"11001101",	-- 0x1073
		"00101011",	-- 0x1074
		"00001100",	-- 0x1075
		"11011010",	-- 0x1076
		"11110001",	-- 0x1077
		"00010000",	-- 0x1078
		"00100010",	-- 0x1079
		"01010101",	-- 0x107A
		"11111011",	-- 0x107B
		"10101111",	-- 0x107C
		"10111110",	-- 0x107D
		"11001010",	-- 0x107E
		"11110111",	-- 0x107F
		"00010000",	-- 0x1080
		"00111110",	-- 0x1081
		"11100101",	-- 0x1082
		"10111110",	-- 0x1083
		"00101000",	-- 0x1084
		"01001011",	-- 0x1085
		"11011101",	-- 0x1086
		"00101010",	-- 0x1087
		"01010101",	-- 0x1088
		"11111011",	-- 0x1089
		"11011101",	-- 0x108A
		"01111110",	-- 0x108B
		"00001011",	-- 0x108C
		"11111110",	-- 0x108D
		"00001111",	-- 0x108E
		"00101000",	-- 0x108F
		"01000000",	-- 0x1090
		"11001011",	-- 0x1091
		"01100111",	-- 0x1092
		"00100000",	-- 0x1093
		"00111100",	-- 0x1094
		"11011101",	-- 0x1095
		"00110110",	-- 0x1096
		"00001011",	-- 0x1097
		"00000000",	-- 0x1098
		"11101101",	-- 0x1099
		"01011011",	-- 0x109A
		"01010101",	-- 0x109B
		"11111011",	-- 0x109C
		"11111101",	-- 0x109D
		"11100101",	-- 0x109E
		"11100001",	-- 0x109F
		"11001101",	-- 0x10A0
		"11000010",	-- 0x10A1
		"00001010",	-- 0x10A2
		"11111110",	-- 0x10A3
		"00000000",	-- 0x10A4
		"00100000",	-- 0x10A5
		"00101010",	-- 0x10A6
		"11011101",	-- 0x10A7
		"01111110",	-- 0x10A8
		"00011011",	-- 0x10A9
		"11111101",	-- 0x10AA
		"01110111",	-- 0x10AB
		"00010001",	-- 0x10AC
		"11011101",	-- 0x10AD
		"01111110",	-- 0x10AE
		"00011010",	-- 0x10AF
		"11111101",	-- 0x10B0
		"01110111",	-- 0x10B1
		"00010000",	-- 0x10B2
		"11011101",	-- 0x10B3
		"01111110",	-- 0x10B4
		"00011100",	-- 0x10B5
		"11111101",	-- 0x10B6
		"01110111",	-- 0x10B7
		"00001100",	-- 0x10B8
		"11011101",	-- 0x10B9
		"01111110",	-- 0x10BA
		"00011101",	-- 0x10BB
		"11111101",	-- 0x10BC
		"01110111",	-- 0x10BD
		"00001101",	-- 0x10BE
		"11011101",	-- 0x10BF
		"01111110",	-- 0x10C0
		"00011110",	-- 0x10C1
		"11111101",	-- 0x10C2
		"01110111",	-- 0x10C3
		"00001110",	-- 0x10C4
		"11011101",	-- 0x10C5
		"01111110",	-- 0x10C6
		"00011111",	-- 0x10C7
		"11111101",	-- 0x10C8
		"01110111",	-- 0x10C9
		"00001111",	-- 0x10CA
		"11111101",	-- 0x10CB
		"00110110",	-- 0x10CC
		"00010010",	-- 0x10CD
		"00000001",	-- 0x10CE
		"00011000",	-- 0x10CF
		"00100110",	-- 0x10D0
		"00000001",	-- 0x10D1
		"00100000",	-- 0x10D2
		"00000000",	-- 0x10D3
		"00101010",	-- 0x10D4
		"01010101",	-- 0x10D5
		"11111011",	-- 0x10D6
		"00001001",	-- 0x10D7
		"00100010",	-- 0x10D8
		"01010101",	-- 0x10D9
		"11111011",	-- 0x10DA
		"11101101",	-- 0x10DB
		"01001011",	-- 0x10DC
		"01011011",	-- 0x10DD
		"11111011",	-- 0x10DE
		"10100111",	-- 0x10DF
		"11101101",	-- 0x10E0
		"01000010",	-- 0x10E1
		"11000010",	-- 0x10E2
		"01111001",	-- 0x10E3
		"00010000",	-- 0x10E4
		"00100001",	-- 0x10E5
		"01010111",	-- 0x10E6
		"11111011",	-- 0x10E7
		"00110100",	-- 0x10E8
		"11000011",	-- 0x10E9
		"01101000",	-- 0x10EA
		"00010000",	-- 0x10EB
		"00100001",	-- 0x10EC
		"11111101",	-- 0x10ED
		"00010000",	-- 0x10EE
		"00011000",	-- 0x10EF
		"00000011",	-- 0x10F0
		"00100001",	-- 0x10F1
		"00011110",	-- 0x10F2
		"00010001",	-- 0x10F3
		"11001101",	-- 0x10F4
		"01101001",	-- 0x10F5
		"00001011",	-- 0x10F6
		"11011101",	-- 0x10F7
		"11100001",	-- 0x10F8
		"11010001",	-- 0x10F9
		"11000001",	-- 0x10FA
		"11110001",	-- 0x10FB
		"11001001",	-- 0x10FC
		"01000110",	-- 0x10FD
		"01000001",	-- 0x10FE
		"01010100",	-- 0x10FF
		"01000001",	-- 0x1100
		"01001100",	-- 0x1101
		"00101000",	-- 0x1102
		"01000110",	-- 0x1103
		"01001111",	-- 0x1104
		"01010000",	-- 0x1105
		"01000101",	-- 0x1106
		"01001110",	-- 0x1107
		"00101001",	-- 0x1108
		"00111010",	-- 0x1109
		"00100000",	-- 0x110A
		"01001110",	-- 0x110B
		"01101111",	-- 0x110C
		"00100000",	-- 0x110D
		"01100100",	-- 0x110E
		"01101001",	-- 0x110F
		"01110011",	-- 0x1110
		"01101011",	-- 0x1111
		"00100000",	-- 0x1112
		"01101101",	-- 0x1113
		"01101111",	-- 0x1114
		"01110101",	-- 0x1115
		"01101110",	-- 0x1116
		"01110100",	-- 0x1117
		"01100101",	-- 0x1118
		"01100100",	-- 0x1119
		"00100001",	-- 0x111A
		"00001101",	-- 0x111B
		"00001010",	-- 0x111C
		"00000000",	-- 0x111D
		"01000110",	-- 0x111E
		"01000001",	-- 0x111F
		"01010100",	-- 0x1120
		"01000001",	-- 0x1121
		"01001100",	-- 0x1122
		"00101000",	-- 0x1123
		"01000110",	-- 0x1124
		"01001111",	-- 0x1125
		"01010000",	-- 0x1126
		"01000101",	-- 0x1127
		"01001110",	-- 0x1128
		"00101001",	-- 0x1129
		"00111010",	-- 0x112A
		"00100000",	-- 0x112B
		"01000011",	-- 0x112C
		"01101111",	-- 0x112D
		"01110101",	-- 0x112E
		"01101100",	-- 0x112F
		"01100100",	-- 0x1130
		"00100000",	-- 0x1131
		"01101110",	-- 0x1132
		"01101111",	-- 0x1133
		"01110100",	-- 0x1134
		"00100000",	-- 0x1135
		"01110010",	-- 0x1136
		"01100101",	-- 0x1137
		"01100001",	-- 0x1138
		"01100100",	-- 0x1139
		"00100000",	-- 0x113A
		"01100100",	-- 0x113B
		"01101001",	-- 0x113C
		"01110010",	-- 0x113D
		"01100101",	-- 0x113E
		"01100011",	-- 0x113F
		"01110100",	-- 0x1140
		"01101111",	-- 0x1141
		"01110010",	-- 0x1142
		"01111001",	-- 0x1143
		"00100000",	-- 0x1144
		"01110011",	-- 0x1145
		"01100101",	-- 0x1146
		"01100011",	-- 0x1147
		"01110100",	-- 0x1148
		"01101111",	-- 0x1149
		"01110010",	-- 0x114A
		"00100001",	-- 0x114B
		"00001101",	-- 0x114C
		"00001010",	-- 0x114D
		"00000000",	-- 0x114E
		"11110101",	-- 0x114F
		"11100101",	-- 0x1150
		"11011001",	-- 0x1151
		"11000101",	-- 0x1152
		"11010101",	-- 0x1153
		"11100101",	-- 0x1154
		"00000001",	-- 0x1155
		"00000000",	-- 0x1156
		"00000000",	-- 0x1157
		"01010000",	-- 0x1158
		"01011001",	-- 0x1159
		"11011001",	-- 0x115A
		"00000001",	-- 0x115B
		"00000010",	-- 0x115C
		"00000000",	-- 0x115D
		"11101101",	-- 0x115E
		"01000010",	-- 0x115F
		"01000100",	-- 0x1160
		"01001101",	-- 0x1161
		"00111010",	-- 0x1162
		"11100101",	-- 0x1163
		"11111101",	-- 0x1164
		"00010110",	-- 0x1165
		"00000000",	-- 0x1166
		"01011111",	-- 0x1167
		"11001101",	-- 0x1168
		"01010100",	-- 0x1169
		"00001101",	-- 0x116A
		"11101101",	-- 0x116B
		"01011011",	-- 0x116C
		"11111100",	-- 0x116D
		"11111101",	-- 0x116E
		"11011001",	-- 0x116F
		"11101101",	-- 0x1170
		"01011011",	-- 0x1171
		"11111110",	-- 0x1172
		"11111101",	-- 0x1173
		"11011001",	-- 0x1174
		"11001101",	-- 0x1175
		"01001110",	-- 0x1176
		"00001101",	-- 0x1177
		"11011001",	-- 0x1178
		"11100101",	-- 0x1179
		"11011001",	-- 0x117A
		"11000001",	-- 0x117B
		"01010100",	-- 0x117C
		"01011101",	-- 0x117D
		"11011001",	-- 0x117E
		"11100001",	-- 0x117F
		"11010001",	-- 0x1180
		"11000001",	-- 0x1181
		"11011001",	-- 0x1182
		"11100001",	-- 0x1183
		"11110001",	-- 0x1184
		"11001001",	-- 0x1185
		"11110101",	-- 0x1186
		"11000101",	-- 0x1187
		"11010101",	-- 0x1188
		"11100101",	-- 0x1189
		"11011101",	-- 0x118A
		"11100101",	-- 0x118B
		"00100001",	-- 0x118C
		"11011100",	-- 0x118D
		"11111101",	-- 0x118E
		"01111110",	-- 0x118F
		"11111110",	-- 0x1190
		"00000000",	-- 0x1191
		"11001010",	-- 0x1192
		"01011001",	-- 0x1193
		"00010010",	-- 0x1194
		"11011101",	-- 0x1195
		"00100001",	-- 0x1196
		"01101101",	-- 0x1197
		"11111011",	-- 0x1198
		"11011101",	-- 0x1199
		"00110110",	-- 0x119A
		"00001000",	-- 0x119B
		"00101110",	-- 0x119C
		"11011101",	-- 0x119D
		"00110110",	-- 0x119E
		"00001100",	-- 0x119F
		"00000000",	-- 0x11A0
		"00100001",	-- 0x11A1
		"10001001",	-- 0x11A2
		"00010010",	-- 0x11A3
		"11001101",	-- 0x11A4
		"01101001",	-- 0x11A5
		"00001011",	-- 0x11A6
		"00100001",	-- 0x11A7
		"00000000",	-- 0x11A8
		"11111110",	-- 0x11A9
		"00000001",	-- 0x11AA
		"00000000",	-- 0x11AB
		"00000010",	-- 0x11AC
		"00001001",	-- 0x11AD
		"00100010",	-- 0x11AE
		"01010001",	-- 0x11AF
		"11111011",	-- 0x11B0
		"00101010",	-- 0x11B1
		"11111000",	-- 0x11B2
		"11111101",	-- 0x11B3
		"00100010",	-- 0x11B4
		"01001101",	-- 0x11B5
		"11111011",	-- 0x11B6
		"00101010",	-- 0x11B7
		"11111010",	-- 0x11B8
		"11111101",	-- 0x11B9
		"00100010",	-- 0x11BA
		"01001111",	-- 0x11BB
		"11111011",	-- 0x11BC
		"11101101",	-- 0x11BD
		"01001011",	-- 0x11BE
		"01001111",	-- 0x11BF
		"11111011",	-- 0x11C0
		"11101101",	-- 0x11C1
		"01011011",	-- 0x11C2
		"01001101",	-- 0x11C3
		"11111011",	-- 0x11C4
		"00100001",	-- 0x11C5
		"00000000",	-- 0x11C6
		"11111110",	-- 0x11C7
		"11001101",	-- 0x11C8
		"00101011",	-- 0x11C9
		"00001100",	-- 0x11CA
		"11011010",	-- 0x11CB
		"01010100",	-- 0x11CC
		"00010010",	-- 0x11CD
		"10101111",	-- 0x11CE
		"10111110",	-- 0x11CF
		"11001010",	-- 0x11D0
		"01011111",	-- 0x11D1
		"00010010",	-- 0x11D2
		"00111110",	-- 0x11D3
		"11100101",	-- 0x11D4
		"10111110",	-- 0x11D5
		"00101000",	-- 0x11D6
		"01100111",	-- 0x11D7
		"00100010",	-- 0x11D8
		"01010011",	-- 0x11D9
		"11111011",	-- 0x11DA
		"11011101",	-- 0x11DB
		"00101010",	-- 0x11DC
		"01010011",	-- 0x11DD
		"11111011",	-- 0x11DE
		"11011101",	-- 0x11DF
		"01111110",	-- 0x11E0
		"00001011",	-- 0x11E1
		"11111110",	-- 0x11E2
		"00001111",	-- 0x11E3
		"00101000",	-- 0x11E4
		"01011001",	-- 0x11E5
		"00010001",	-- 0x11E6
		"01101101",	-- 0x11E7
		"11111011",	-- 0x11E8
		"00000001",	-- 0x11E9
		"00001000",	-- 0x11EA
		"00000000",	-- 0x11EB
		"11101101",	-- 0x11EC
		"10110000",	-- 0x11ED
		"00010011",	-- 0x11EE
		"00000001",	-- 0x11EF
		"00000011",	-- 0x11F0
		"00000000",	-- 0x11F1
		"11101101",	-- 0x11F2
		"10110000",	-- 0x11F3
		"00100001",	-- 0x11F4
		"01101101",	-- 0x11F5
		"11111011",	-- 0x11F6
		"11001101",	-- 0x11F7
		"01101001",	-- 0x11F8
		"00001011",	-- 0x11F9
		"00100001",	-- 0x11FA
		"01011110",	-- 0x11FB
		"00010011",	-- 0x11FC
		"11001011",	-- 0x11FD
		"01100111",	-- 0x11FE
		"00101000",	-- 0x11FF
		"00000011",	-- 0x1200
		"00100001",	-- 0x1201
		"01011000",	-- 0x1202
		"00010011",	-- 0x1203
		"11001101",	-- 0x1204
		"01101001",	-- 0x1205
		"00001011",	-- 0x1206
		"11011101",	-- 0x1207
		"01100110",	-- 0x1208
		"00011111",	-- 0x1209
		"11011101",	-- 0x120A
		"01101110",	-- 0x120B
		"00011110",	-- 0x120C
		"11001101",	-- 0x120D
		"01010110",	-- 0x120E
		"00001011",	-- 0x120F
		"11011101",	-- 0x1210
		"01100110",	-- 0x1211
		"00011101",	-- 0x1212
		"11011101",	-- 0x1213
		"01101110",	-- 0x1214
		"00011100",	-- 0x1215
		"11001101",	-- 0x1216
		"01010110",	-- 0x1217
		"00001011",	-- 0x1218
		"00111110",	-- 0x1219
		"00001001",	-- 0x121A
		"11001101",	-- 0x121B
		"01100011",	-- 0x121C
		"00001011",	-- 0x121D
		"11011101",	-- 0x121E
		"01100110",	-- 0x121F
		"00011011",	-- 0x1220
		"11011101",	-- 0x1221
		"01101110",	-- 0x1222
		"00011010",	-- 0x1223
		"00000001",	-- 0x1224
		"00000000",	-- 0x1225
		"00000000",	-- 0x1226
		"10100111",	-- 0x1227
		"11101101",	-- 0x1228
		"01000010",	-- 0x1229
		"00101000",	-- 0x122A
		"00001101",	-- 0x122B
		"11001101",	-- 0x122C
		"01001111",	-- 0x122D
		"00010001",	-- 0x122E
		"01100000",	-- 0x122F
		"01101001",	-- 0x1230
		"11001101",	-- 0x1231
		"01010110",	-- 0x1232
		"00001011",	-- 0x1233
		"01100010",	-- 0x1234
		"01101011",	-- 0x1235
		"11001101",	-- 0x1236
		"01010110",	-- 0x1237
		"00001011",	-- 0x1238
		"11001101",	-- 0x1239
		"11010100",	-- 0x123A
		"00001010",	-- 0x123B
		"00101010",	-- 0x123C
		"01010011",	-- 0x123D
		"11111011",	-- 0x123E
		"00000001",	-- 0x123F
		"00100000",	-- 0x1240
		"00000000",	-- 0x1241
		"00001001",	-- 0x1242
		"11101101",	-- 0x1243
		"01001011",	-- 0x1244
		"01010001",	-- 0x1245
		"11111011",	-- 0x1246
		"10100111",	-- 0x1247
		"11101101",	-- 0x1248
		"01000010",	-- 0x1249
		"11000010",	-- 0x124A
		"11001110",	-- 0x124B
		"00010001",	-- 0x124C
		"00100001",	-- 0x124D
		"01001101",	-- 0x124E
		"11111011",	-- 0x124F
		"00110100",	-- 0x1250
		"11000011",	-- 0x1251
		"10111101",	-- 0x1252
		"00010001",	-- 0x1253
		"00100001",	-- 0x1254
		"00100110",	-- 0x1255
		"00010011",	-- 0x1256
		"00011000",	-- 0x1257
		"00000011",	-- 0x1258
		"00100001",	-- 0x1259
		"01100110",	-- 0x125A
		"00010010",	-- 0x125B
		"11001101",	-- 0x125C
		"01101001",	-- 0x125D
		"00001011",	-- 0x125E
		"11011101",	-- 0x125F
		"11100001",	-- 0x1260
		"11100001",	-- 0x1261
		"11010001",	-- 0x1262
		"11000001",	-- 0x1263
		"11110001",	-- 0x1264
		"11001001",	-- 0x1265
		"01000110",	-- 0x1266
		"01000001",	-- 0x1267
		"01010100",	-- 0x1268
		"01000001",	-- 0x1269
		"01001100",	-- 0x126A
		"00101000",	-- 0x126B
		"01000100",	-- 0x126C
		"01001001",	-- 0x126D
		"01010010",	-- 0x126E
		"01001100",	-- 0x126F
		"01001001",	-- 0x1270
		"01010011",	-- 0x1271
		"01010100",	-- 0x1272
		"00101001",	-- 0x1273
		"00111010",	-- 0x1274
		"00100000",	-- 0x1275
		"01001110",	-- 0x1276
		"01101111",	-- 0x1277
		"00100000",	-- 0x1278
		"01100100",	-- 0x1279
		"01101001",	-- 0x127A
		"01110011",	-- 0x127B
		"01101011",	-- 0x127C
		"00100000",	-- 0x127D
		"01101101",	-- 0x127E
		"01101111",	-- 0x127F
		"01110101",	-- 0x1280
		"01101110",	-- 0x1281
		"01110100",	-- 0x1282
		"01100101",	-- 0x1283
		"01100100",	-- 0x1284
		"00100001",	-- 0x1285
		"00001101",	-- 0x1286
		"00001010",	-- 0x1287
		"00000000",	-- 0x1288
		"01000100",	-- 0x1289
		"01101001",	-- 0x128A
		"01110010",	-- 0x128B
		"01100101",	-- 0x128C
		"01100011",	-- 0x128D
		"01110100",	-- 0x128E
		"01101111",	-- 0x128F
		"01110010",	-- 0x1290
		"01111001",	-- 0x1291
		"00100000",	-- 0x1292
		"01100011",	-- 0x1293
		"01101111",	-- 0x1294
		"01101110",	-- 0x1295
		"01110100",	-- 0x1296
		"01100101",	-- 0x1297
		"01101110",	-- 0x1298
		"01110100",	-- 0x1299
		"01110011",	-- 0x129A
		"00111010",	-- 0x129B
		"00001101",	-- 0x129C
		"00001010",	-- 0x129D
		"00101101",	-- 0x129E
		"00101101",	-- 0x129F
		"00101101",	-- 0x12A0
		"00101101",	-- 0x12A1
		"00101101",	-- 0x12A2
		"00101101",	-- 0x12A3
		"00101101",	-- 0x12A4
		"00101101",	-- 0x12A5
		"00101101",	-- 0x12A6
		"00101101",	-- 0x12A7
		"00101101",	-- 0x12A8
		"00101101",	-- 0x12A9
		"00101101",	-- 0x12AA
		"00101101",	-- 0x12AB
		"00101101",	-- 0x12AC
		"00101101",	-- 0x12AD
		"00101101",	-- 0x12AE
		"00101101",	-- 0x12AF
		"00101101",	-- 0x12B0
		"00101101",	-- 0x12B1
		"00101101",	-- 0x12B2
		"00101101",	-- 0x12B3
		"00101101",	-- 0x12B4
		"00101101",	-- 0x12B5
		"00101101",	-- 0x12B6
		"00101101",	-- 0x12B7
		"00101101",	-- 0x12B8
		"00101101",	-- 0x12B9
		"00101101",	-- 0x12BA
		"00101101",	-- 0x12BB
		"00101101",	-- 0x12BC
		"00101101",	-- 0x12BD
		"00101101",	-- 0x12BE
		"00101101",	-- 0x12BF
		"00101101",	-- 0x12C0
		"00101101",	-- 0x12C1
		"00101101",	-- 0x12C2
		"00101101",	-- 0x12C3
		"00101101",	-- 0x12C4
		"00101101",	-- 0x12C5
		"00101101",	-- 0x12C6
		"00101101",	-- 0x12C7
		"00101101",	-- 0x12C8
		"00001101",	-- 0x12C9
		"00001010",	-- 0x12CA
		"01000110",	-- 0x12CB
		"01001001",	-- 0x12CC
		"01001100",	-- 0x12CD
		"01000101",	-- 0x12CE
		"01001110",	-- 0x12CF
		"01000001",	-- 0x12D0
		"01001101",	-- 0x12D1
		"01000101",	-- 0x12D2
		"00101110",	-- 0x12D3
		"01000101",	-- 0x12D4
		"01011000",	-- 0x12D5
		"01010100",	-- 0x12D6
		"00100000",	-- 0x12D7
		"00100000",	-- 0x12D8
		"01000100",	-- 0x12D9
		"01001001",	-- 0x12DA
		"01010010",	-- 0x12DB
		"00111111",	-- 0x12DC
		"00100000",	-- 0x12DD
		"00100000",	-- 0x12DE
		"00100000",	-- 0x12DF
		"01010011",	-- 0x12E0
		"01001001",	-- 0x12E1
		"01011010",	-- 0x12E2
		"01000101",	-- 0x12E3
		"00100000",	-- 0x12E4
		"00101000",	-- 0x12E5
		"01000010",	-- 0x12E6
		"01011001",	-- 0x12E7
		"01010100",	-- 0x12E8
		"01000101",	-- 0x12E9
		"01010011",	-- 0x12EA
		"00101001",	-- 0x12EB
		"00100000",	-- 0x12EC
		"00100000",	-- 0x12ED
		"00110001",	-- 0x12EE
		"01010011",	-- 0x12EF
		"01010100",	-- 0x12F0
		"00100000",	-- 0x12F1
		"01010011",	-- 0x12F2
		"01000101",	-- 0x12F3
		"01000011",	-- 0x12F4
		"01010100",	-- 0x12F5
		"00001101",	-- 0x12F6
		"00001010",	-- 0x12F7
		"00101101",	-- 0x12F8
		"00101101",	-- 0x12F9
		"00101101",	-- 0x12FA
		"00101101",	-- 0x12FB
		"00101101",	-- 0x12FC
		"00101101",	-- 0x12FD
		"00101101",	-- 0x12FE
		"00101101",	-- 0x12FF
		"00101101",	-- 0x1300
		"00101101",	-- 0x1301
		"00101101",	-- 0x1302
		"00101101",	-- 0x1303
		"00101101",	-- 0x1304
		"00101101",	-- 0x1305
		"00101101",	-- 0x1306
		"00101101",	-- 0x1307
		"00101101",	-- 0x1308
		"00101101",	-- 0x1309
		"00101101",	-- 0x130A
		"00101101",	-- 0x130B
		"00101101",	-- 0x130C
		"00101101",	-- 0x130D
		"00101101",	-- 0x130E
		"00101101",	-- 0x130F
		"00101101",	-- 0x1310
		"00101101",	-- 0x1311
		"00101101",	-- 0x1312
		"00101101",	-- 0x1313
		"00101101",	-- 0x1314
		"00101101",	-- 0x1315
		"00101101",	-- 0x1316
		"00101101",	-- 0x1317
		"00101101",	-- 0x1318
		"00101101",	-- 0x1319
		"00101101",	-- 0x131A
		"00101101",	-- 0x131B
		"00101101",	-- 0x131C
		"00101101",	-- 0x131D
		"00101101",	-- 0x131E
		"00101101",	-- 0x131F
		"00101101",	-- 0x1320
		"00101101",	-- 0x1321
		"00101101",	-- 0x1322
		"00001101",	-- 0x1323
		"00001010",	-- 0x1324
		"00000000",	-- 0x1325
		"01000110",	-- 0x1326
		"01000001",	-- 0x1327
		"01010100",	-- 0x1328
		"01000001",	-- 0x1329
		"01001100",	-- 0x132A
		"00101000",	-- 0x132B
		"01000100",	-- 0x132C
		"01001001",	-- 0x132D
		"01010010",	-- 0x132E
		"01001100",	-- 0x132F
		"01001001",	-- 0x1330
		"01010011",	-- 0x1331
		"01010100",	-- 0x1332
		"00101001",	-- 0x1333
		"00111010",	-- 0x1334
		"00100000",	-- 0x1335
		"01000011",	-- 0x1336
		"01101111",	-- 0x1337
		"01110101",	-- 0x1338
		"01101100",	-- 0x1339
		"01100100",	-- 0x133A
		"00100000",	-- 0x133B
		"01101110",	-- 0x133C
		"01101111",	-- 0x133D
		"01110100",	-- 0x133E
		"00100000",	-- 0x133F
		"01110010",	-- 0x1340
		"01100101",	-- 0x1341
		"01100001",	-- 0x1342
		"01100100",	-- 0x1343
		"00100000",	-- 0x1344
		"01100100",	-- 0x1345
		"01101001",	-- 0x1346
		"01110010",	-- 0x1347
		"01100101",	-- 0x1348
		"01100011",	-- 0x1349
		"01110100",	-- 0x134A
		"01101111",	-- 0x134B
		"01110010",	-- 0x134C
		"01111001",	-- 0x134D
		"00100000",	-- 0x134E
		"01110011",	-- 0x134F
		"01100101",	-- 0x1350
		"01100011",	-- 0x1351
		"01110100",	-- 0x1352
		"01101111",	-- 0x1353
		"01110010",	-- 0x1354
		"00001101",	-- 0x1355
		"00001010",	-- 0x1356
		"00000000",	-- 0x1357
		"00001001",	-- 0x1358
		"01000100",	-- 0x1359
		"01001001",	-- 0x135A
		"01010010",	-- 0x135B
		"00001001",	-- 0x135C
		"00000000",	-- 0x135D
		"00001001",	-- 0x135E
		"00001001",	-- 0x135F
		"00000000",	-- 0x1360
		"11110101",	-- 0x1361
		"11000101",	-- 0x1362
		"11010101",	-- 0x1363
		"11100101",	-- 0x1364
		"11011101",	-- 0x1365
		"11100101",	-- 0x1366
		"00100001",	-- 0x1367
		"00000000",	-- 0x1368
		"11111110",	-- 0x1369
		"00000001",	-- 0x136A
		"00000000",	-- 0x136B
		"00000000",	-- 0x136C
		"00010001",	-- 0x136D
		"00000000",	-- 0x136E
		"00000000",	-- 0x136F
		"11001101",	-- 0x1370
		"00101011",	-- 0x1371
		"00001100",	-- 0x1372
		"11011010",	-- 0x1373
		"11011001",	-- 0x1374
		"00010100",	-- 0x1375
		"11011101",	-- 0x1376
		"00100001",	-- 0x1377
		"11111110",	-- 0x1378
		"11111111",	-- 0x1379
		"00111110",	-- 0x137A
		"01010101",	-- 0x137B
		"11011101",	-- 0x137C
		"10111110",	-- 0x137D
		"00000000",	-- 0x137E
		"11000010",	-- 0x137F
		"11011110",	-- 0x1380
		"00010100",	-- 0x1381
		"00111110",	-- 0x1382
		"10101010",	-- 0x1383
		"11011101",	-- 0x1384
		"10111110",	-- 0x1385
		"00000001",	-- 0x1386
		"11000010",	-- 0x1387
		"11011110",	-- 0x1388
		"00010100",	-- 0x1389
		"00000001",	-- 0x138A
		"00001000",	-- 0x138B
		"00000000",	-- 0x138C
		"00100001",	-- 0x138D
		"11000110",	-- 0x138E
		"11111111",	-- 0x138F
		"00010001",	-- 0x1390
		"11101100",	-- 0x1391
		"11111101",	-- 0x1392
		"11101101",	-- 0x1393
		"10110000",	-- 0x1394
		"00100001",	-- 0x1395
		"00000000",	-- 0x1396
		"11111110",	-- 0x1397
		"11101101",	-- 0x1398
		"01011011",	-- 0x1399
		"11101100",	-- 0x139A
		"11111101",	-- 0x139B
		"11101101",	-- 0x139C
		"01001011",	-- 0x139D
		"11101110",	-- 0x139E
		"11111101",	-- 0x139F
		"11001101",	-- 0x13A0
		"00101011",	-- 0x13A1
		"00001100",	-- 0x13A2
		"11011010",	-- 0x13A3
		"11100011",	-- 0x13A4
		"00010100",	-- 0x13A5
		"00000001",	-- 0x13A6
		"00001000",	-- 0x13A7
		"00000000",	-- 0x13A8
		"00100001",	-- 0x13A9
		"00000011",	-- 0x13AA
		"11111110",	-- 0x13AB
		"00010001",	-- 0x13AC
		"11011100",	-- 0x13AD
		"11111101",	-- 0x13AE
		"11101101",	-- 0x13AF
		"10110000",	-- 0x13B0
		"11011101",	-- 0x13B1
		"00100001",	-- 0x13B2
		"00000000",	-- 0x13B3
		"11111110",	-- 0x13B4
		"00111110",	-- 0x13B5
		"00000010",	-- 0x13B6
		"11011101",	-- 0x13B7
		"10111110",	-- 0x13B8
		"00010000",	-- 0x13B9
		"11000010",	-- 0x13BA
		"11101000",	-- 0x13BB
		"00010100",	-- 0x13BC
		"10101111",	-- 0x13BD
		"11011101",	-- 0x13BE
		"10111110",	-- 0x13BF
		"00001011",	-- 0x13C0
		"11000010",	-- 0x13C1
		"11101101",	-- 0x13C2
		"00010100",	-- 0x13C3
		"00111110",	-- 0x13C4
		"00000010",	-- 0x13C5
		"11011101",	-- 0x13C6
		"10111110",	-- 0x13C7
		"00001100",	-- 0x13C8
		"11000010",	-- 0x13C9
		"11101101",	-- 0x13CA
		"00010100",	-- 0x13CB
		"00111010",	-- 0x13CC
		"00001101",	-- 0x13CD
		"11111110",	-- 0x13CE
		"00110010",	-- 0x13CF
		"11100101",	-- 0x13D0
		"11111101",	-- 0x13D1
		"11101101",	-- 0x13D2
		"01001011",	-- 0x13D3
		"00001110",	-- 0x13D4
		"11111110",	-- 0x13D5
		"11101101",	-- 0x13D6
		"01000011",	-- 0x13D7
		"11100110",	-- 0x13D8
		"11111101",	-- 0x13D9
		"11101101",	-- 0x13DA
		"01001011",	-- 0x13DB
		"00010110",	-- 0x13DC
		"11111110",	-- 0x13DD
		"11101101",	-- 0x13DE
		"01000011",	-- 0x13DF
		"11101000",	-- 0x13E0
		"11111101",	-- 0x13E1
		"11101101",	-- 0x13E2
		"01001011",	-- 0x13E3
		"00010001",	-- 0x13E4
		"11111110",	-- 0x13E5
		"11101101",	-- 0x13E6
		"01000011",	-- 0x13E7
		"11101010",	-- 0x13E8
		"11111101",	-- 0x13E9
		"00101010",	-- 0x13EA
		"11101100",	-- 0x13EB
		"11111101",	-- 0x13EC
		"11101101",	-- 0x13ED
		"01001011",	-- 0x13EE
		"11100110",	-- 0x13EF
		"11111101",	-- 0x13F0
		"00001001",	-- 0x13F1
		"00100010",	-- 0x13F2
		"11110100",	-- 0x13F3
		"11111101",	-- 0x13F4
		"00101010",	-- 0x13F5
		"11101110",	-- 0x13F6
		"11111101",	-- 0x13F7
		"00000001",	-- 0x13F8
		"00000000",	-- 0x13F9
		"00000000",	-- 0x13FA
		"11101101",	-- 0x13FB
		"01001010",	-- 0x13FC
		"00100010",	-- 0x13FD
		"11110110",	-- 0x13FE
		"11111101",	-- 0x13FF
		"00101010",	-- 0x1400
		"11101000",	-- 0x1401
		"11111101",	-- 0x1402
		"00101001",	-- 0x1403
		"01000100",	-- 0x1404
		"01001101",	-- 0x1405
		"00101010",	-- 0x1406
		"11110100",	-- 0x1407
		"11111101",	-- 0x1408
		"00001001",	-- 0x1409
		"00100010",	-- 0x140A
		"11111000",	-- 0x140B
		"11111101",	-- 0x140C
		"00101010",	-- 0x140D
		"11110110",	-- 0x140E
		"11111101",	-- 0x140F
		"00000001",	-- 0x1410
		"00000000",	-- 0x1411
		"00000000",	-- 0x1412
		"11101101",	-- 0x1413
		"01001010",	-- 0x1414
		"00100010",	-- 0x1415
		"11111010",	-- 0x1416
		"11111101",	-- 0x1417
		"11101101",	-- 0x1418
		"01001011",	-- 0x1419
		"11101010",	-- 0x141A
		"11111101",	-- 0x141B
		"11001011",	-- 0x141C
		"00101000",	-- 0x141D
		"11001011",	-- 0x141E
		"00011001",	-- 0x141F
		"11001011",	-- 0x1420
		"00101000",	-- 0x1421
		"11001011",	-- 0x1422
		"00011001",	-- 0x1423
		"11001011",	-- 0x1424
		"00101000",	-- 0x1425
		"11001011",	-- 0x1426
		"00011001",	-- 0x1427
		"11001011",	-- 0x1428
		"00101000",	-- 0x1429
		"11001011",	-- 0x142A
		"00011001",	-- 0x142B
		"00101010",	-- 0x142C
		"11111000",	-- 0x142D
		"11111101",	-- 0x142E
		"00001001",	-- 0x142F
		"00100010",	-- 0x1430
		"11111100",	-- 0x1431
		"11111101",	-- 0x1432
		"00101010",	-- 0x1433
		"11111010",	-- 0x1434
		"11111101",	-- 0x1435
		"00000001",	-- 0x1436
		"00000000",	-- 0x1437
		"00000000",	-- 0x1438
		"11101101",	-- 0x1439
		"01001010",	-- 0x143A
		"00100010",	-- 0x143B
		"11111110",	-- 0x143C
		"11111101",	-- 0x143D
		"00100001",	-- 0x143E
		"11011001",	-- 0x143F
		"00010101",	-- 0x1440
		"11001101",	-- 0x1441
		"01101001",	-- 0x1442
		"00001011",	-- 0x1443
		"00100001",	-- 0x1444
		"11011100",	-- 0x1445
		"11111101",	-- 0x1446
		"11001101",	-- 0x1447
		"01101001",	-- 0x1448
		"00001011",	-- 0x1449
		"00100001",	-- 0x144A
		"11100100",	-- 0x144B
		"00010101",	-- 0x144C
		"11001101",	-- 0x144D
		"01101001",	-- 0x144E
		"00001011",	-- 0x144F
		"00111010",	-- 0x1450
		"11100101",	-- 0x1451
		"11111101",	-- 0x1452
		"11001101",	-- 0x1453
		"00110101",	-- 0x1454
		"00001011",	-- 0x1455
		"00100001",	-- 0x1456
		"11110000",	-- 0x1457
		"00010101",	-- 0x1458
		"11001101",	-- 0x1459
		"01101001",	-- 0x145A
		"00001011",	-- 0x145B
		"00101010",	-- 0x145C
		"11100110",	-- 0x145D
		"11111101",	-- 0x145E
		"11001101",	-- 0x145F
		"01010110",	-- 0x1460
		"00001011",	-- 0x1461
		"00100001",	-- 0x1462
		"11111100",	-- 0x1463
		"00010101",	-- 0x1464
		"11001101",	-- 0x1465
		"01101001",	-- 0x1466
		"00001011",	-- 0x1467
		"00101010",	-- 0x1468
		"11101000",	-- 0x1469
		"11111101",	-- 0x146A
		"11001101",	-- 0x146B
		"01010110",	-- 0x146C
		"00001011",	-- 0x146D
		"00100001",	-- 0x146E
		"00001000",	-- 0x146F
		"00010110",	-- 0x1470
		"11001101",	-- 0x1471
		"01101001",	-- 0x1472
		"00001011",	-- 0x1473
		"00101010",	-- 0x1474
		"11101010",	-- 0x1475
		"11111101",	-- 0x1476
		"11001101",	-- 0x1477
		"01010110",	-- 0x1478
		"00001011",	-- 0x1479
		"00100001",	-- 0x147A
		"00010101",	-- 0x147B
		"00010110",	-- 0x147C
		"11001101",	-- 0x147D
		"01101001",	-- 0x147E
		"00001011",	-- 0x147F
		"00101010",	-- 0x1480
		"11110010",	-- 0x1481
		"11111101",	-- 0x1482
		"11001101",	-- 0x1483
		"01010110",	-- 0x1484
		"00001011",	-- 0x1485
		"00101010",	-- 0x1486
		"11110000",	-- 0x1487
		"11111101",	-- 0x1488
		"11001101",	-- 0x1489
		"01010110",	-- 0x148A
		"00001011",	-- 0x148B
		"00100001",	-- 0x148C
		"00100000",	-- 0x148D
		"00010110",	-- 0x148E
		"11001101",	-- 0x148F
		"01101001",	-- 0x1490
		"00001011",	-- 0x1491
		"00101010",	-- 0x1492
		"11101110",	-- 0x1493
		"11111101",	-- 0x1494
		"11001101",	-- 0x1495
		"01010110",	-- 0x1496
		"00001011",	-- 0x1497
		"00101010",	-- 0x1498
		"11101100",	-- 0x1499
		"11111101",	-- 0x149A
		"11001101",	-- 0x149B
		"01010110",	-- 0x149C
		"00001011",	-- 0x149D
		"00100001",	-- 0x149E
		"00101100",	-- 0x149F
		"00010110",	-- 0x14A0
		"11001101",	-- 0x14A1
		"01101001",	-- 0x14A2
		"00001011",	-- 0x14A3
		"00101010",	-- 0x14A4
		"11110110",	-- 0x14A5
		"11111101",	-- 0x14A6
		"11001101",	-- 0x14A7
		"01010110",	-- 0x14A8
		"00001011",	-- 0x14A9
		"00101010",	-- 0x14AA
		"11110100",	-- 0x14AB
		"11111101",	-- 0x14AC
		"11001101",	-- 0x14AD
		"01010110",	-- 0x14AE
		"00001011",	-- 0x14AF
		"00100001",	-- 0x14B0
		"00111011",	-- 0x14B1
		"00010110",	-- 0x14B2
		"11001101",	-- 0x14B3
		"01101001",	-- 0x14B4
		"00001011",	-- 0x14B5
		"00101010",	-- 0x14B6
		"11111010",	-- 0x14B7
		"11111101",	-- 0x14B8
		"11001101",	-- 0x14B9
		"01010110",	-- 0x14BA
		"00001011",	-- 0x14BB
		"00101010",	-- 0x14BC
		"11111000",	-- 0x14BD
		"11111101",	-- 0x14BE
		"11001101",	-- 0x14BF
		"01010110",	-- 0x14C0
		"00001011",	-- 0x14C1
		"00100001",	-- 0x14C2
		"01001010",	-- 0x14C3
		"00010110",	-- 0x14C4
		"11001101",	-- 0x14C5
		"01101001",	-- 0x14C6
		"00001011",	-- 0x14C7
		"00101010",	-- 0x14C8
		"11111110",	-- 0x14C9
		"11111101",	-- 0x14CA
		"11001101",	-- 0x14CB
		"01010110",	-- 0x14CC
		"00001011",	-- 0x14CD
		"00101010",	-- 0x14CE
		"11111100",	-- 0x14CF
		"11111101",	-- 0x14D0
		"11001101",	-- 0x14D1
		"01010110",	-- 0x14D2
		"00001011",	-- 0x14D3
		"11001101",	-- 0x14D4
		"11010100",	-- 0x14D5
		"00001010",	-- 0x14D6
		"00011000",	-- 0x14D7
		"00011010",	-- 0x14D8
		"00100001",	-- 0x14D9
		"11111010",	-- 0x14DA
		"00010100",	-- 0x14DB
		"00011000",	-- 0x14DC
		"00010010",	-- 0x14DD
		"00100001",	-- 0x14DE
		"00100001",	-- 0x14DF
		"00010101",	-- 0x14E0
		"00011000",	-- 0x14E1
		"00001101",	-- 0x14E2
		"00100001",	-- 0x14E3
		"01000001",	-- 0x14E4
		"00010101",	-- 0x14E5
		"00011000",	-- 0x14E6
		"00001000",	-- 0x14E7
		"00100001",	-- 0x14E8
		"01111000",	-- 0x14E9
		"00010101",	-- 0x14EA
		"00011000",	-- 0x14EB
		"00000011",	-- 0x14EC
		"00100001",	-- 0x14ED
		"10100101",	-- 0x14EE
		"00010101",	-- 0x14EF
		"11001101",	-- 0x14F0
		"01101001",	-- 0x14F1
		"00001011",	-- 0x14F2
		"11011101",	-- 0x14F3
		"11100001",	-- 0x14F4
		"11100001",	-- 0x14F5
		"11010001",	-- 0x14F6
		"11000001",	-- 0x14F7
		"11110001",	-- 0x14F8
		"11001001",	-- 0x14F9
		"01000110",	-- 0x14FA
		"01000001",	-- 0x14FB
		"01010100",	-- 0x14FC
		"01000001",	-- 0x14FD
		"01001100",	-- 0x14FE
		"00101000",	-- 0x14FF
		"01000110",	-- 0x1500
		"01000001",	-- 0x1501
		"01010100",	-- 0x1502
		"01001101",	-- 0x1503
		"01001111",	-- 0x1504
		"01010101",	-- 0x1505
		"01001110",	-- 0x1506
		"01010100",	-- 0x1507
		"00101001",	-- 0x1508
		"00111010",	-- 0x1509
		"00100000",	-- 0x150A
		"01000011",	-- 0x150B
		"01101111",	-- 0x150C
		"01110101",	-- 0x150D
		"01101100",	-- 0x150E
		"01100100",	-- 0x150F
		"00100000",	-- 0x1510
		"01101110",	-- 0x1511
		"01101111",	-- 0x1512
		"01110100",	-- 0x1513
		"00100000",	-- 0x1514
		"01110010",	-- 0x1515
		"01100101",	-- 0x1516
		"01100001",	-- 0x1517
		"01100100",	-- 0x1518
		"00100000",	-- 0x1519
		"01001101",	-- 0x151A
		"01000010",	-- 0x151B
		"01010010",	-- 0x151C
		"00100001",	-- 0x151D
		"00001101",	-- 0x151E
		"00001010",	-- 0x151F
		"00000000",	-- 0x1520
		"01000110",	-- 0x1521
		"01000001",	-- 0x1522
		"01010100",	-- 0x1523
		"01000001",	-- 0x1524
		"01001100",	-- 0x1525
		"00101000",	-- 0x1526
		"01000110",	-- 0x1527
		"01000001",	-- 0x1528
		"01010100",	-- 0x1529
		"01001101",	-- 0x152A
		"01001111",	-- 0x152B
		"01010101",	-- 0x152C
		"01001110",	-- 0x152D
		"01010100",	-- 0x152E
		"00101001",	-- 0x152F
		"00111010",	-- 0x1530
		"00100000",	-- 0x1531
		"01001001",	-- 0x1532
		"01101100",	-- 0x1533
		"01101100",	-- 0x1534
		"01100101",	-- 0x1535
		"01100111",	-- 0x1536
		"01100001",	-- 0x1537
		"01101100",	-- 0x1538
		"00100000",	-- 0x1539
		"01001101",	-- 0x153A
		"01000010",	-- 0x153B
		"01010010",	-- 0x153C
		"00100001",	-- 0x153D
		"00001101",	-- 0x153E
		"00001010",	-- 0x153F
		"00000000",	-- 0x1540
		"01000110",	-- 0x1541
		"01000001",	-- 0x1542
		"01010100",	-- 0x1543
		"01000001",	-- 0x1544
		"01001100",	-- 0x1545
		"00101000",	-- 0x1546
		"01000110",	-- 0x1547
		"01000001",	-- 0x1548
		"01010100",	-- 0x1549
		"01001101",	-- 0x154A
		"01001111",	-- 0x154B
		"01010101",	-- 0x154C
		"01001110",	-- 0x154D
		"01010100",	-- 0x154E
		"00101001",	-- 0x154F
		"00111010",	-- 0x1550
		"00100000",	-- 0x1551
		"01000011",	-- 0x1552
		"01101111",	-- 0x1553
		"01110101",	-- 0x1554
		"01101100",	-- 0x1555
		"01100100",	-- 0x1556
		"00100000",	-- 0x1557
		"01101110",	-- 0x1558
		"01101111",	-- 0x1559
		"01110100",	-- 0x155A
		"00100000",	-- 0x155B
		"01110010",	-- 0x155C
		"01100101",	-- 0x155D
		"01100001",	-- 0x155E
		"01100100",	-- 0x155F
		"00100000",	-- 0x1560
		"01110000",	-- 0x1561
		"01100001",	-- 0x1562
		"01110010",	-- 0x1563
		"01110100",	-- 0x1564
		"01101001",	-- 0x1565
		"01110100",	-- 0x1566
		"01101001",	-- 0x1567
		"01101111",	-- 0x1568
		"01101110",	-- 0x1569
		"00100000",	-- 0x156A
		"01100010",	-- 0x156B
		"01101111",	-- 0x156C
		"01101111",	-- 0x156D
		"01110100",	-- 0x156E
		"00100000",	-- 0x156F
		"01100010",	-- 0x1570
		"01101100",	-- 0x1571
		"01101111",	-- 0x1572
		"01100011",	-- 0x1573
		"01101011",	-- 0x1574
		"00001101",	-- 0x1575
		"00001010",	-- 0x1576
		"00000000",	-- 0x1577
		"01000110",	-- 0x1578
		"01000001",	-- 0x1579
		"01010100",	-- 0x157A
		"01000001",	-- 0x157B
		"01001100",	-- 0x157C
		"00101000",	-- 0x157D
		"01000110",	-- 0x157E
		"01000001",	-- 0x157F
		"01010100",	-- 0x1580
		"01001101",	-- 0x1581
		"01001111",	-- 0x1582
		"01010101",	-- 0x1583
		"01001110",	-- 0x1584
		"01010100",	-- 0x1585
		"00101001",	-- 0x1586
		"00111010",	-- 0x1587
		"00100000",	-- 0x1588
		"01000110",	-- 0x1589
		"01000001",	-- 0x158A
		"01010100",	-- 0x158B
		"00100000",	-- 0x158C
		"01101110",	-- 0x158D
		"01110101",	-- 0x158E
		"01101101",	-- 0x158F
		"01100010",	-- 0x1590
		"01100101",	-- 0x1591
		"01110010",	-- 0x1592
		"00100000",	-- 0x1593
		"01101110",	-- 0x1594
		"01101111",	-- 0x1595
		"01110100",	-- 0x1596
		"00100000",	-- 0x1597
		"01100101",	-- 0x1598
		"01110001",	-- 0x1599
		"01110101",	-- 0x159A
		"01100001",	-- 0x159B
		"01101100",	-- 0x159C
		"00100000",	-- 0x159D
		"01110100",	-- 0x159E
		"01110111",	-- 0x159F
		"01101111",	-- 0x15A0
		"00100001",	-- 0x15A1
		"00001101",	-- 0x15A2
		"00001010",	-- 0x15A3
		"00000000",	-- 0x15A4
		"01000110",	-- 0x15A5
		"01000001",	-- 0x15A6
		"01010100",	-- 0x15A7
		"01000001",	-- 0x15A8
		"01001100",	-- 0x15A9
		"00101000",	-- 0x15AA
		"01000110",	-- 0x15AB
		"01000001",	-- 0x15AC
		"01010100",	-- 0x15AD
		"01001101",	-- 0x15AE
		"01001111",	-- 0x15AF
		"01010101",	-- 0x15B0
		"01001110",	-- 0x15B1
		"01010100",	-- 0x15B2
		"00101001",	-- 0x15B3
		"00111010",	-- 0x15B4
		"00100000",	-- 0x15B5
		"01010011",	-- 0x15B6
		"01100101",	-- 0x15B7
		"01100011",	-- 0x15B8
		"01110100",	-- 0x15B9
		"01101111",	-- 0x15BA
		"01110010",	-- 0x15BB
		"00100000",	-- 0x15BC
		"01110011",	-- 0x15BD
		"01101001",	-- 0x15BE
		"01111010",	-- 0x15BF
		"01100101",	-- 0x15C0
		"00100000",	-- 0x15C1
		"01101110",	-- 0x15C2
		"01101111",	-- 0x15C3
		"01110100",	-- 0x15C4
		"00100000",	-- 0x15C5
		"01100101",	-- 0x15C6
		"01110001",	-- 0x15C7
		"01110101",	-- 0x15C8
		"01100001",	-- 0x15C9
		"01101100",	-- 0x15CA
		"00100000",	-- 0x15CB
		"00110101",	-- 0x15CC
		"00110001",	-- 0x15CD
		"00110010",	-- 0x15CE
		"00100000",	-- 0x15CF
		"01100010",	-- 0x15D0
		"01111001",	-- 0x15D1
		"01110100",	-- 0x15D2
		"01100101",	-- 0x15D3
		"01110011",	-- 0x15D4
		"00100001",	-- 0x15D5
		"00001101",	-- 0x15D6
		"00001010",	-- 0x15D7
		"00000000",	-- 0x15D8
		"00001001",	-- 0x15D9
		"01000110",	-- 0x15DA
		"01000001",	-- 0x15DB
		"01010100",	-- 0x15DC
		"01001110",	-- 0x15DD
		"01000001",	-- 0x15DE
		"01001101",	-- 0x15DF
		"01000101",	-- 0x15E0
		"00111010",	-- 0x15E1
		"00001001",	-- 0x15E2
		"00000000",	-- 0x15E3
		"00001101",	-- 0x15E4
		"00001010",	-- 0x15E5
		"00001001",	-- 0x15E6
		"01000011",	-- 0x15E7
		"01001100",	-- 0x15E8
		"01010101",	-- 0x15E9
		"01010011",	-- 0x15EA
		"01001001",	-- 0x15EB
		"01011010",	-- 0x15EC
		"00111010",	-- 0x15ED
		"00001001",	-- 0x15EE
		"00000000",	-- 0x15EF
		"00001101",	-- 0x15F0
		"00001010",	-- 0x15F1
		"00001001",	-- 0x15F2
		"01010010",	-- 0x15F3
		"01000101",	-- 0x15F4
		"01010011",	-- 0x15F5
		"01010011",	-- 0x15F6
		"01000101",	-- 0x15F7
		"01000011",	-- 0x15F8
		"00111010",	-- 0x15F9
		"00001001",	-- 0x15FA
		"00000000",	-- 0x15FB
		"00001101",	-- 0x15FC
		"00001010",	-- 0x15FD
		"00001001",	-- 0x15FE
		"01000110",	-- 0x15FF
		"01000001",	-- 0x1600
		"01010100",	-- 0x1601
		"01010011",	-- 0x1602
		"01000101",	-- 0x1603
		"01000011",	-- 0x1604
		"00111010",	-- 0x1605
		"00001001",	-- 0x1606
		"00000000",	-- 0x1607
		"00001101",	-- 0x1608
		"00001010",	-- 0x1609
		"00001001",	-- 0x160A
		"01010010",	-- 0x160B
		"01001111",	-- 0x160C
		"01001111",	-- 0x160D
		"01010100",	-- 0x160E
		"01001100",	-- 0x160F
		"01000101",	-- 0x1610
		"01001110",	-- 0x1611
		"00111010",	-- 0x1612
		"00001001",	-- 0x1613
		"00000000",	-- 0x1614
		"00001101",	-- 0x1615
		"00001010",	-- 0x1616
		"00001001",	-- 0x1617
		"01010000",	-- 0x1618
		"01010011",	-- 0x1619
		"01001001",	-- 0x161A
		"01011010",	-- 0x161B
		"00111010",	-- 0x161C
		"00001001",	-- 0x161D
		"00001001",	-- 0x161E
		"00000000",	-- 0x161F
		"00001101",	-- 0x1620
		"00001010",	-- 0x1621
		"00001001",	-- 0x1622
		"01010000",	-- 0x1623
		"01010011",	-- 0x1624
		"01010100",	-- 0x1625
		"01000001",	-- 0x1626
		"01010010",	-- 0x1627
		"01010100",	-- 0x1628
		"00111010",	-- 0x1629
		"00001001",	-- 0x162A
		"00000000",	-- 0x162B
		"00001101",	-- 0x162C
		"00001010",	-- 0x162D
		"00001001",	-- 0x162E
		"01000110",	-- 0x162F
		"01000001",	-- 0x1630
		"01010100",	-- 0x1631
		"00110001",	-- 0x1632
		"01010011",	-- 0x1633
		"01010100",	-- 0x1634
		"01000001",	-- 0x1635
		"01010010",	-- 0x1636
		"01010100",	-- 0x1637
		"00111010",	-- 0x1638
		"00001001",	-- 0x1639
		"00000000",	-- 0x163A
		"00001101",	-- 0x163B
		"00001010",	-- 0x163C
		"00001001",	-- 0x163D
		"01010010",	-- 0x163E
		"01001111",	-- 0x163F
		"01001111",	-- 0x1640
		"01010100",	-- 0x1641
		"01010011",	-- 0x1642
		"01010100",	-- 0x1643
		"01000001",	-- 0x1644
		"01010010",	-- 0x1645
		"01010100",	-- 0x1646
		"00111010",	-- 0x1647
		"00001001",	-- 0x1648
		"00000000",	-- 0x1649
		"00001101",	-- 0x164A
		"00001010",	-- 0x164B
		"00001001",	-- 0x164C
		"01000100",	-- 0x164D
		"01000001",	-- 0x164E
		"01010100",	-- 0x164F
		"01000001",	-- 0x1650
		"01010011",	-- 0x1651
		"01010100",	-- 0x1652
		"01000001",	-- 0x1653
		"01010010",	-- 0x1654
		"01010100",	-- 0x1655
		"00111010",	-- 0x1656
		"00001001",	-- 0x1657
		"00000000",	-- 0x1658
		"11110101",	-- 0x1659
		"11100101",	-- 0x165A
		"10101111",	-- 0x165B
		"00100001",	-- 0x165C
		"11011100",	-- 0x165D
		"11111101",	-- 0x165E
		"01110111",	-- 0x165F
		"11100001",	-- 0x1660
		"11110001",	-- 0x1661
		"11001001",	-- 0x1662
		"01010100",	-- 0x1663
		"01001000",	-- 0x1664
		"01000101",	-- 0x1665
		"00100000",	-- 0x1666
		"01001101",	-- 0x1667
		"01001111",	-- 0x1668
		"01001110",	-- 0x1669
		"01001001",	-- 0x166A
		"01010100",	-- 0x166B
		"01001111",	-- 0x166C
		"01010010",	-- 0x166D
		"00100000",	-- 0x166E
		"01000101",	-- 0x166F
		"01001110",	-- 0x1670
		"01000100",	-- 0x1671
		"01010011",	-- 0x1672
		"00100000",	-- 0x1673
		"01001000",	-- 0x1674
		"01000101",	-- 0x1675
		"01010010",	-- 0x1676
		"01000101",	-- 0x1677
		"00101110",	-- 0x1678
		"00101110",	-- 0x1679
		"00101110",	-- 0x167A
		"00000000",	-- 0x167B
		"--------",	-- 0x167C
		"--------",	-- 0x167D
		"--------",	-- 0x167E
		"--------",	-- 0x167F
		"--------",	-- 0x1680
		"--------",	-- 0x1681
		"--------",	-- 0x1682
		"--------",	-- 0x1683
		"--------",	-- 0x1684
		"--------",	-- 0x1685
		"--------",	-- 0x1686
		"--------",	-- 0x1687
		"--------",	-- 0x1688
		"--------",	-- 0x1689
		"--------",	-- 0x168A
		"--------",	-- 0x168B
		"--------",	-- 0x168C
		"--------",	-- 0x168D
		"--------",	-- 0x168E
		"--------",	-- 0x168F
		"--------",	-- 0x1690
		"--------",	-- 0x1691
		"--------",	-- 0x1692
		"--------",	-- 0x1693
		"--------",	-- 0x1694
		"--------",	-- 0x1695
		"--------",	-- 0x1696
		"--------",	-- 0x1697
		"--------",	-- 0x1698
		"--------",	-- 0x1699
		"--------",	-- 0x169A
		"--------",	-- 0x169B
		"--------",	-- 0x169C
		"--------",	-- 0x169D
		"--------",	-- 0x169E
		"--------",	-- 0x169F
		"--------",	-- 0x16A0
		"--------",	-- 0x16A1
		"--------",	-- 0x16A2
		"--------",	-- 0x16A3
		"--------",	-- 0x16A4
		"--------",	-- 0x16A5
		"--------",	-- 0x16A6
		"--------",	-- 0x16A7
		"--------",	-- 0x16A8
		"--------",	-- 0x16A9
		"--------",	-- 0x16AA
		"--------",	-- 0x16AB
		"--------",	-- 0x16AC
		"--------",	-- 0x16AD
		"--------",	-- 0x16AE
		"--------",	-- 0x16AF
		"--------",	-- 0x16B0
		"--------",	-- 0x16B1
		"--------",	-- 0x16B2
		"--------",	-- 0x16B3
		"--------",	-- 0x16B4
		"--------",	-- 0x16B5
		"--------",	-- 0x16B6
		"--------",	-- 0x16B7
		"--------",	-- 0x16B8
		"--------",	-- 0x16B9
		"--------",	-- 0x16BA
		"--------",	-- 0x16BB
		"--------",	-- 0x16BC
		"--------",	-- 0x16BD
		"--------",	-- 0x16BE
		"--------",	-- 0x16BF
		"--------",	-- 0x16C0
		"--------",	-- 0x16C1
		"--------",	-- 0x16C2
		"--------",	-- 0x16C3
		"--------",	-- 0x16C4
		"--------",	-- 0x16C5
		"--------",	-- 0x16C6
		"--------",	-- 0x16C7
		"--------",	-- 0x16C8
		"--------",	-- 0x16C9
		"--------",	-- 0x16CA
		"--------",	-- 0x16CB
		"--------",	-- 0x16CC
		"--------",	-- 0x16CD
		"--------",	-- 0x16CE
		"--------",	-- 0x16CF
		"--------",	-- 0x16D0
		"--------",	-- 0x16D1
		"--------",	-- 0x16D2
		"--------",	-- 0x16D3
		"--------",	-- 0x16D4
		"--------",	-- 0x16D5
		"--------",	-- 0x16D6
		"--------",	-- 0x16D7
		"--------",	-- 0x16D8
		"--------",	-- 0x16D9
		"--------",	-- 0x16DA
		"--------",	-- 0x16DB
		"--------",	-- 0x16DC
		"--------",	-- 0x16DD
		"--------",	-- 0x16DE
		"--------",	-- 0x16DF
		"--------",	-- 0x16E0
		"--------",	-- 0x16E1
		"--------",	-- 0x16E2
		"--------",	-- 0x16E3
		"--------",	-- 0x16E4
		"--------",	-- 0x16E5
		"--------",	-- 0x16E6
		"--------",	-- 0x16E7
		"--------",	-- 0x16E8
		"--------",	-- 0x16E9
		"--------",	-- 0x16EA
		"--------",	-- 0x16EB
		"--------",	-- 0x16EC
		"--------",	-- 0x16ED
		"--------",	-- 0x16EE
		"--------",	-- 0x16EF
		"--------",	-- 0x16F0
		"--------",	-- 0x16F1
		"--------",	-- 0x16F2
		"--------",	-- 0x16F3
		"--------",	-- 0x16F4
		"--------",	-- 0x16F5
		"--------",	-- 0x16F6
		"--------",	-- 0x16F7
		"--------",	-- 0x16F8
		"--------",	-- 0x16F9
		"--------",	-- 0x16FA
		"--------",	-- 0x16FB
		"--------",	-- 0x16FC
		"--------",	-- 0x16FD
		"--------",	-- 0x16FE
		"--------",	-- 0x16FF
		"--------",	-- 0x1700
		"--------",	-- 0x1701
		"--------",	-- 0x1702
		"--------",	-- 0x1703
		"--------",	-- 0x1704
		"--------",	-- 0x1705
		"--------",	-- 0x1706
		"--------",	-- 0x1707
		"--------",	-- 0x1708
		"--------",	-- 0x1709
		"--------",	-- 0x170A
		"--------",	-- 0x170B
		"--------",	-- 0x170C
		"--------",	-- 0x170D
		"--------",	-- 0x170E
		"--------",	-- 0x170F
		"--------",	-- 0x1710
		"--------",	-- 0x1711
		"--------",	-- 0x1712
		"--------",	-- 0x1713
		"--------",	-- 0x1714
		"--------",	-- 0x1715
		"--------",	-- 0x1716
		"--------",	-- 0x1717
		"--------",	-- 0x1718
		"--------",	-- 0x1719
		"--------",	-- 0x171A
		"--------",	-- 0x171B
		"--------",	-- 0x171C
		"--------",	-- 0x171D
		"--------",	-- 0x171E
		"--------",	-- 0x171F
		"--------",	-- 0x1720
		"--------",	-- 0x1721
		"--------",	-- 0x1722
		"--------",	-- 0x1723
		"--------",	-- 0x1724
		"--------",	-- 0x1725
		"--------",	-- 0x1726
		"--------",	-- 0x1727
		"--------",	-- 0x1728
		"--------",	-- 0x1729
		"--------",	-- 0x172A
		"--------",	-- 0x172B
		"--------",	-- 0x172C
		"--------",	-- 0x172D
		"--------",	-- 0x172E
		"--------",	-- 0x172F
		"--------",	-- 0x1730
		"--------",	-- 0x1731
		"--------",	-- 0x1732
		"--------",	-- 0x1733
		"--------",	-- 0x1734
		"--------",	-- 0x1735
		"--------",	-- 0x1736
		"--------",	-- 0x1737
		"--------",	-- 0x1738
		"--------",	-- 0x1739
		"--------",	-- 0x173A
		"--------",	-- 0x173B
		"--------",	-- 0x173C
		"--------",	-- 0x173D
		"--------",	-- 0x173E
		"--------",	-- 0x173F
		"--------",	-- 0x1740
		"--------",	-- 0x1741
		"--------",	-- 0x1742
		"--------",	-- 0x1743
		"--------",	-- 0x1744
		"--------",	-- 0x1745
		"--------",	-- 0x1746
		"--------",	-- 0x1747
		"--------",	-- 0x1748
		"--------",	-- 0x1749
		"--------",	-- 0x174A
		"--------",	-- 0x174B
		"--------",	-- 0x174C
		"--------",	-- 0x174D
		"--------",	-- 0x174E
		"--------",	-- 0x174F
		"--------",	-- 0x1750
		"--------",	-- 0x1751
		"--------",	-- 0x1752
		"--------",	-- 0x1753
		"--------",	-- 0x1754
		"--------",	-- 0x1755
		"--------",	-- 0x1756
		"--------",	-- 0x1757
		"--------",	-- 0x1758
		"--------",	-- 0x1759
		"--------",	-- 0x175A
		"--------",	-- 0x175B
		"--------",	-- 0x175C
		"--------",	-- 0x175D
		"--------",	-- 0x175E
		"--------",	-- 0x175F
		"--------",	-- 0x1760
		"--------",	-- 0x1761
		"--------",	-- 0x1762
		"--------",	-- 0x1763
		"--------",	-- 0x1764
		"--------",	-- 0x1765
		"--------",	-- 0x1766
		"--------",	-- 0x1767
		"--------",	-- 0x1768
		"--------",	-- 0x1769
		"--------",	-- 0x176A
		"--------",	-- 0x176B
		"--------",	-- 0x176C
		"--------",	-- 0x176D
		"--------",	-- 0x176E
		"--------",	-- 0x176F
		"--------",	-- 0x1770
		"--------",	-- 0x1771
		"--------",	-- 0x1772
		"--------",	-- 0x1773
		"--------",	-- 0x1774
		"--------",	-- 0x1775
		"--------",	-- 0x1776
		"--------",	-- 0x1777
		"--------",	-- 0x1778
		"--------",	-- 0x1779
		"--------",	-- 0x177A
		"--------",	-- 0x177B
		"--------",	-- 0x177C
		"--------",	-- 0x177D
		"--------",	-- 0x177E
		"--------",	-- 0x177F
		"--------",	-- 0x1780
		"--------",	-- 0x1781
		"--------",	-- 0x1782
		"--------",	-- 0x1783
		"--------",	-- 0x1784
		"--------",	-- 0x1785
		"--------",	-- 0x1786
		"--------",	-- 0x1787
		"--------",	-- 0x1788
		"--------",	-- 0x1789
		"--------",	-- 0x178A
		"--------",	-- 0x178B
		"--------",	-- 0x178C
		"--------",	-- 0x178D
		"--------",	-- 0x178E
		"--------",	-- 0x178F
		"--------",	-- 0x1790
		"--------",	-- 0x1791
		"--------",	-- 0x1792
		"--------",	-- 0x1793
		"--------",	-- 0x1794
		"--------",	-- 0x1795
		"--------",	-- 0x1796
		"--------",	-- 0x1797
		"--------",	-- 0x1798
		"--------",	-- 0x1799
		"--------",	-- 0x179A
		"--------",	-- 0x179B
		"--------",	-- 0x179C
		"--------",	-- 0x179D
		"--------",	-- 0x179E
		"--------",	-- 0x179F
		"--------",	-- 0x17A0
		"--------",	-- 0x17A1
		"--------",	-- 0x17A2
		"--------",	-- 0x17A3
		"--------",	-- 0x17A4
		"--------",	-- 0x17A5
		"--------",	-- 0x17A6
		"--------",	-- 0x17A7
		"--------",	-- 0x17A8
		"--------",	-- 0x17A9
		"--------",	-- 0x17AA
		"--------",	-- 0x17AB
		"--------",	-- 0x17AC
		"--------",	-- 0x17AD
		"--------",	-- 0x17AE
		"--------",	-- 0x17AF
		"--------",	-- 0x17B0
		"--------",	-- 0x17B1
		"--------",	-- 0x17B2
		"--------",	-- 0x17B3
		"--------",	-- 0x17B4
		"--------",	-- 0x17B5
		"--------",	-- 0x17B6
		"--------",	-- 0x17B7
		"--------",	-- 0x17B8
		"--------",	-- 0x17B9
		"--------",	-- 0x17BA
		"--------",	-- 0x17BB
		"--------",	-- 0x17BC
		"--------",	-- 0x17BD
		"--------",	-- 0x17BE
		"--------",	-- 0x17BF
		"--------",	-- 0x17C0
		"--------",	-- 0x17C1
		"--------",	-- 0x17C2
		"--------",	-- 0x17C3
		"--------",	-- 0x17C4
		"--------",	-- 0x17C5
		"--------",	-- 0x17C6
		"--------",	-- 0x17C7
		"--------",	-- 0x17C8
		"--------",	-- 0x17C9
		"--------",	-- 0x17CA
		"--------",	-- 0x17CB
		"--------",	-- 0x17CC
		"--------",	-- 0x17CD
		"--------",	-- 0x17CE
		"--------",	-- 0x17CF
		"--------",	-- 0x17D0
		"--------",	-- 0x17D1
		"--------",	-- 0x17D2
		"--------",	-- 0x17D3
		"--------",	-- 0x17D4
		"--------",	-- 0x17D5
		"--------",	-- 0x17D6
		"--------",	-- 0x17D7
		"--------",	-- 0x17D8
		"--------",	-- 0x17D9
		"--------",	-- 0x17DA
		"--------",	-- 0x17DB
		"--------",	-- 0x17DC
		"--------",	-- 0x17DD
		"--------",	-- 0x17DE
		"--------",	-- 0x17DF
		"--------",	-- 0x17E0
		"--------",	-- 0x17E1
		"--------",	-- 0x17E2
		"--------",	-- 0x17E3
		"--------",	-- 0x17E4
		"--------",	-- 0x17E5
		"--------",	-- 0x17E6
		"--------",	-- 0x17E7
		"--------",	-- 0x17E8
		"--------",	-- 0x17E9
		"--------",	-- 0x17EA
		"--------",	-- 0x17EB
		"--------",	-- 0x17EC
		"--------",	-- 0x17ED
		"--------",	-- 0x17EE
		"--------",	-- 0x17EF
		"--------",	-- 0x17F0
		"--------",	-- 0x17F1
		"--------",	-- 0x17F2
		"--------",	-- 0x17F3
		"--------",	-- 0x17F4
		"--------",	-- 0x17F5
		"--------",	-- 0x17F6
		"--------",	-- 0x17F7
		"--------",	-- 0x17F8
		"--------",	-- 0x17F9
		"--------",	-- 0x17FA
		"--------",	-- 0x17FB
		"--------",	-- 0x17FC
		"--------",	-- 0x17FD
		"--------",	-- 0x17FE
		"--------",	-- 0x17FF
		"--------",	-- 0x1800
		"--------",	-- 0x1801
		"--------",	-- 0x1802
		"--------",	-- 0x1803
		"--------",	-- 0x1804
		"--------",	-- 0x1805
		"--------",	-- 0x1806
		"--------",	-- 0x1807
		"--------",	-- 0x1808
		"--------",	-- 0x1809
		"--------",	-- 0x180A
		"--------",	-- 0x180B
		"--------",	-- 0x180C
		"--------",	-- 0x180D
		"--------",	-- 0x180E
		"--------",	-- 0x180F
		"--------",	-- 0x1810
		"--------",	-- 0x1811
		"--------",	-- 0x1812
		"--------",	-- 0x1813
		"--------",	-- 0x1814
		"--------",	-- 0x1815
		"--------",	-- 0x1816
		"--------",	-- 0x1817
		"--------",	-- 0x1818
		"--------",	-- 0x1819
		"--------",	-- 0x181A
		"--------",	-- 0x181B
		"--------",	-- 0x181C
		"--------",	-- 0x181D
		"--------",	-- 0x181E
		"--------",	-- 0x181F
		"--------",	-- 0x1820
		"--------",	-- 0x1821
		"--------",	-- 0x1822
		"--------",	-- 0x1823
		"--------",	-- 0x1824
		"--------",	-- 0x1825
		"--------",	-- 0x1826
		"--------",	-- 0x1827
		"--------",	-- 0x1828
		"--------",	-- 0x1829
		"--------",	-- 0x182A
		"--------",	-- 0x182B
		"--------",	-- 0x182C
		"--------",	-- 0x182D
		"--------",	-- 0x182E
		"--------",	-- 0x182F
		"--------",	-- 0x1830
		"--------",	-- 0x1831
		"--------",	-- 0x1832
		"--------",	-- 0x1833
		"--------",	-- 0x1834
		"--------",	-- 0x1835
		"--------",	-- 0x1836
		"--------",	-- 0x1837
		"--------",	-- 0x1838
		"--------",	-- 0x1839
		"--------",	-- 0x183A
		"--------",	-- 0x183B
		"--------",	-- 0x183C
		"--------",	-- 0x183D
		"--------",	-- 0x183E
		"--------",	-- 0x183F
		"--------",	-- 0x1840
		"--------",	-- 0x1841
		"--------",	-- 0x1842
		"--------",	-- 0x1843
		"--------",	-- 0x1844
		"--------",	-- 0x1845
		"--------",	-- 0x1846
		"--------",	-- 0x1847
		"--------",	-- 0x1848
		"--------",	-- 0x1849
		"--------",	-- 0x184A
		"--------",	-- 0x184B
		"--------",	-- 0x184C
		"--------",	-- 0x184D
		"--------",	-- 0x184E
		"--------",	-- 0x184F
		"--------",	-- 0x1850
		"--------",	-- 0x1851
		"--------",	-- 0x1852
		"--------",	-- 0x1853
		"--------",	-- 0x1854
		"--------",	-- 0x1855
		"--------",	-- 0x1856
		"--------",	-- 0x1857
		"--------",	-- 0x1858
		"--------",	-- 0x1859
		"--------",	-- 0x185A
		"--------",	-- 0x185B
		"--------",	-- 0x185C
		"--------",	-- 0x185D
		"--------",	-- 0x185E
		"--------",	-- 0x185F
		"--------",	-- 0x1860
		"--------",	-- 0x1861
		"--------",	-- 0x1862
		"--------",	-- 0x1863
		"--------",	-- 0x1864
		"--------",	-- 0x1865
		"--------",	-- 0x1866
		"--------",	-- 0x1867
		"--------",	-- 0x1868
		"--------",	-- 0x1869
		"--------",	-- 0x186A
		"--------",	-- 0x186B
		"--------",	-- 0x186C
		"--------",	-- 0x186D
		"--------",	-- 0x186E
		"--------",	-- 0x186F
		"--------",	-- 0x1870
		"--------",	-- 0x1871
		"--------",	-- 0x1872
		"--------",	-- 0x1873
		"--------",	-- 0x1874
		"--------",	-- 0x1875
		"--------",	-- 0x1876
		"--------",	-- 0x1877
		"--------",	-- 0x1878
		"--------",	-- 0x1879
		"--------",	-- 0x187A
		"--------",	-- 0x187B
		"--------",	-- 0x187C
		"--------",	-- 0x187D
		"--------",	-- 0x187E
		"--------",	-- 0x187F
		"--------",	-- 0x1880
		"--------",	-- 0x1881
		"--------",	-- 0x1882
		"--------",	-- 0x1883
		"--------",	-- 0x1884
		"--------",	-- 0x1885
		"--------",	-- 0x1886
		"--------",	-- 0x1887
		"--------",	-- 0x1888
		"--------",	-- 0x1889
		"--------",	-- 0x188A
		"--------",	-- 0x188B
		"--------",	-- 0x188C
		"--------",	-- 0x188D
		"--------",	-- 0x188E
		"--------",	-- 0x188F
		"--------",	-- 0x1890
		"--------",	-- 0x1891
		"--------",	-- 0x1892
		"--------",	-- 0x1893
		"--------",	-- 0x1894
		"--------",	-- 0x1895
		"--------",	-- 0x1896
		"--------",	-- 0x1897
		"--------",	-- 0x1898
		"--------",	-- 0x1899
		"--------",	-- 0x189A
		"--------",	-- 0x189B
		"--------",	-- 0x189C
		"--------",	-- 0x189D
		"--------",	-- 0x189E
		"--------",	-- 0x189F
		"--------",	-- 0x18A0
		"--------",	-- 0x18A1
		"--------",	-- 0x18A2
		"--------",	-- 0x18A3
		"--------",	-- 0x18A4
		"--------",	-- 0x18A5
		"--------",	-- 0x18A6
		"--------",	-- 0x18A7
		"--------",	-- 0x18A8
		"--------",	-- 0x18A9
		"--------",	-- 0x18AA
		"--------",	-- 0x18AB
		"--------",	-- 0x18AC
		"--------",	-- 0x18AD
		"--------",	-- 0x18AE
		"--------",	-- 0x18AF
		"--------",	-- 0x18B0
		"--------",	-- 0x18B1
		"--------",	-- 0x18B2
		"--------",	-- 0x18B3
		"--------",	-- 0x18B4
		"--------",	-- 0x18B5
		"--------",	-- 0x18B6
		"--------",	-- 0x18B7
		"--------",	-- 0x18B8
		"--------",	-- 0x18B9
		"--------",	-- 0x18BA
		"--------",	-- 0x18BB
		"--------",	-- 0x18BC
		"--------",	-- 0x18BD
		"--------",	-- 0x18BE
		"--------",	-- 0x18BF
		"--------",	-- 0x18C0
		"--------",	-- 0x18C1
		"--------",	-- 0x18C2
		"--------",	-- 0x18C3
		"--------",	-- 0x18C4
		"--------",	-- 0x18C5
		"--------",	-- 0x18C6
		"--------",	-- 0x18C7
		"--------",	-- 0x18C8
		"--------",	-- 0x18C9
		"--------",	-- 0x18CA
		"--------",	-- 0x18CB
		"--------",	-- 0x18CC
		"--------",	-- 0x18CD
		"--------",	-- 0x18CE
		"--------",	-- 0x18CF
		"--------",	-- 0x18D0
		"--------",	-- 0x18D1
		"--------",	-- 0x18D2
		"--------",	-- 0x18D3
		"--------",	-- 0x18D4
		"--------",	-- 0x18D5
		"--------",	-- 0x18D6
		"--------",	-- 0x18D7
		"--------",	-- 0x18D8
		"--------",	-- 0x18D9
		"--------",	-- 0x18DA
		"--------",	-- 0x18DB
		"--------",	-- 0x18DC
		"--------",	-- 0x18DD
		"--------",	-- 0x18DE
		"--------",	-- 0x18DF
		"--------",	-- 0x18E0
		"--------",	-- 0x18E1
		"--------",	-- 0x18E2
		"--------",	-- 0x18E3
		"--------",	-- 0x18E4
		"--------",	-- 0x18E5
		"--------",	-- 0x18E6
		"--------",	-- 0x18E7
		"--------",	-- 0x18E8
		"--------",	-- 0x18E9
		"--------",	-- 0x18EA
		"--------",	-- 0x18EB
		"--------",	-- 0x18EC
		"--------",	-- 0x18ED
		"--------",	-- 0x18EE
		"--------",	-- 0x18EF
		"--------",	-- 0x18F0
		"--------",	-- 0x18F1
		"--------",	-- 0x18F2
		"--------",	-- 0x18F3
		"--------",	-- 0x18F4
		"--------",	-- 0x18F5
		"--------",	-- 0x18F6
		"--------",	-- 0x18F7
		"--------",	-- 0x18F8
		"--------",	-- 0x18F9
		"--------",	-- 0x18FA
		"--------",	-- 0x18FB
		"--------",	-- 0x18FC
		"--------",	-- 0x18FD
		"--------",	-- 0x18FE
		"--------",	-- 0x18FF
		"--------",	-- 0x1900
		"--------",	-- 0x1901
		"--------",	-- 0x1902
		"--------",	-- 0x1903
		"--------",	-- 0x1904
		"--------",	-- 0x1905
		"--------",	-- 0x1906
		"--------",	-- 0x1907
		"--------",	-- 0x1908
		"--------",	-- 0x1909
		"--------",	-- 0x190A
		"--------",	-- 0x190B
		"--------",	-- 0x190C
		"--------",	-- 0x190D
		"--------",	-- 0x190E
		"--------",	-- 0x190F
		"--------",	-- 0x1910
		"--------",	-- 0x1911
		"--------",	-- 0x1912
		"--------",	-- 0x1913
		"--------",	-- 0x1914
		"--------",	-- 0x1915
		"--------",	-- 0x1916
		"--------",	-- 0x1917
		"--------",	-- 0x1918
		"--------",	-- 0x1919
		"--------",	-- 0x191A
		"--------",	-- 0x191B
		"--------",	-- 0x191C
		"--------",	-- 0x191D
		"--------",	-- 0x191E
		"--------",	-- 0x191F
		"--------",	-- 0x1920
		"--------",	-- 0x1921
		"--------",	-- 0x1922
		"--------",	-- 0x1923
		"--------",	-- 0x1924
		"--------",	-- 0x1925
		"--------",	-- 0x1926
		"--------",	-- 0x1927
		"--------",	-- 0x1928
		"--------",	-- 0x1929
		"--------",	-- 0x192A
		"--------",	-- 0x192B
		"--------",	-- 0x192C
		"--------",	-- 0x192D
		"--------",	-- 0x192E
		"--------",	-- 0x192F
		"--------",	-- 0x1930
		"--------",	-- 0x1931
		"--------",	-- 0x1932
		"--------",	-- 0x1933
		"--------",	-- 0x1934
		"--------",	-- 0x1935
		"--------",	-- 0x1936
		"--------",	-- 0x1937
		"--------",	-- 0x1938
		"--------",	-- 0x1939
		"--------",	-- 0x193A
		"--------",	-- 0x193B
		"--------",	-- 0x193C
		"--------",	-- 0x193D
		"--------",	-- 0x193E
		"--------",	-- 0x193F
		"--------",	-- 0x1940
		"--------",	-- 0x1941
		"--------",	-- 0x1942
		"--------",	-- 0x1943
		"--------",	-- 0x1944
		"--------",	-- 0x1945
		"--------",	-- 0x1946
		"--------",	-- 0x1947
		"--------",	-- 0x1948
		"--------",	-- 0x1949
		"--------",	-- 0x194A
		"--------",	-- 0x194B
		"--------",	-- 0x194C
		"--------",	-- 0x194D
		"--------",	-- 0x194E
		"--------",	-- 0x194F
		"--------",	-- 0x1950
		"--------",	-- 0x1951
		"--------",	-- 0x1952
		"--------",	-- 0x1953
		"--------",	-- 0x1954
		"--------",	-- 0x1955
		"--------",	-- 0x1956
		"--------",	-- 0x1957
		"--------",	-- 0x1958
		"--------",	-- 0x1959
		"--------",	-- 0x195A
		"--------",	-- 0x195B
		"--------",	-- 0x195C
		"--------",	-- 0x195D
		"--------",	-- 0x195E
		"--------",	-- 0x195F
		"--------",	-- 0x1960
		"--------",	-- 0x1961
		"--------",	-- 0x1962
		"--------",	-- 0x1963
		"--------",	-- 0x1964
		"--------",	-- 0x1965
		"--------",	-- 0x1966
		"--------",	-- 0x1967
		"--------",	-- 0x1968
		"--------",	-- 0x1969
		"--------",	-- 0x196A
		"--------",	-- 0x196B
		"--------",	-- 0x196C
		"--------",	-- 0x196D
		"--------",	-- 0x196E
		"--------",	-- 0x196F
		"--------",	-- 0x1970
		"--------",	-- 0x1971
		"--------",	-- 0x1972
		"--------",	-- 0x1973
		"--------",	-- 0x1974
		"--------",	-- 0x1975
		"--------",	-- 0x1976
		"--------",	-- 0x1977
		"--------",	-- 0x1978
		"--------",	-- 0x1979
		"--------",	-- 0x197A
		"--------",	-- 0x197B
		"--------",	-- 0x197C
		"--------",	-- 0x197D
		"--------",	-- 0x197E
		"--------",	-- 0x197F
		"--------",	-- 0x1980
		"--------",	-- 0x1981
		"--------",	-- 0x1982
		"--------",	-- 0x1983
		"--------",	-- 0x1984
		"--------",	-- 0x1985
		"--------",	-- 0x1986
		"--------",	-- 0x1987
		"--------",	-- 0x1988
		"--------",	-- 0x1989
		"--------",	-- 0x198A
		"--------",	-- 0x198B
		"--------",	-- 0x198C
		"--------",	-- 0x198D
		"--------",	-- 0x198E
		"--------",	-- 0x198F
		"--------",	-- 0x1990
		"--------",	-- 0x1991
		"--------",	-- 0x1992
		"--------",	-- 0x1993
		"--------",	-- 0x1994
		"--------",	-- 0x1995
		"--------",	-- 0x1996
		"--------",	-- 0x1997
		"--------",	-- 0x1998
		"--------",	-- 0x1999
		"--------",	-- 0x199A
		"--------",	-- 0x199B
		"--------",	-- 0x199C
		"--------",	-- 0x199D
		"--------",	-- 0x199E
		"--------",	-- 0x199F
		"--------",	-- 0x19A0
		"--------",	-- 0x19A1
		"--------",	-- 0x19A2
		"--------",	-- 0x19A3
		"--------",	-- 0x19A4
		"--------",	-- 0x19A5
		"--------",	-- 0x19A6
		"--------",	-- 0x19A7
		"--------",	-- 0x19A8
		"--------",	-- 0x19A9
		"--------",	-- 0x19AA
		"--------",	-- 0x19AB
		"--------",	-- 0x19AC
		"--------",	-- 0x19AD
		"--------",	-- 0x19AE
		"--------",	-- 0x19AF
		"--------",	-- 0x19B0
		"--------",	-- 0x19B1
		"--------",	-- 0x19B2
		"--------",	-- 0x19B3
		"--------",	-- 0x19B4
		"--------",	-- 0x19B5
		"--------",	-- 0x19B6
		"--------",	-- 0x19B7
		"--------",	-- 0x19B8
		"--------",	-- 0x19B9
		"--------",	-- 0x19BA
		"--------",	-- 0x19BB
		"--------",	-- 0x19BC
		"--------",	-- 0x19BD
		"--------",	-- 0x19BE
		"--------",	-- 0x19BF
		"--------",	-- 0x19C0
		"--------",	-- 0x19C1
		"--------",	-- 0x19C2
		"--------",	-- 0x19C3
		"--------",	-- 0x19C4
		"--------",	-- 0x19C5
		"--------",	-- 0x19C6
		"--------",	-- 0x19C7
		"--------",	-- 0x19C8
		"--------",	-- 0x19C9
		"--------",	-- 0x19CA
		"--------",	-- 0x19CB
		"--------",	-- 0x19CC
		"--------",	-- 0x19CD
		"--------",	-- 0x19CE
		"--------",	-- 0x19CF
		"--------",	-- 0x19D0
		"--------",	-- 0x19D1
		"--------",	-- 0x19D2
		"--------",	-- 0x19D3
		"--------",	-- 0x19D4
		"--------",	-- 0x19D5
		"--------",	-- 0x19D6
		"--------",	-- 0x19D7
		"--------",	-- 0x19D8
		"--------",	-- 0x19D9
		"--------",	-- 0x19DA
		"--------",	-- 0x19DB
		"--------",	-- 0x19DC
		"--------",	-- 0x19DD
		"--------",	-- 0x19DE
		"--------",	-- 0x19DF
		"--------",	-- 0x19E0
		"--------",	-- 0x19E1
		"--------",	-- 0x19E2
		"--------",	-- 0x19E3
		"--------",	-- 0x19E4
		"--------",	-- 0x19E5
		"--------",	-- 0x19E6
		"--------",	-- 0x19E7
		"--------",	-- 0x19E8
		"--------",	-- 0x19E9
		"--------",	-- 0x19EA
		"--------",	-- 0x19EB
		"--------",	-- 0x19EC
		"--------",	-- 0x19ED
		"--------",	-- 0x19EE
		"--------",	-- 0x19EF
		"--------",	-- 0x19F0
		"--------",	-- 0x19F1
		"--------",	-- 0x19F2
		"--------",	-- 0x19F3
		"--------",	-- 0x19F4
		"--------",	-- 0x19F5
		"--------",	-- 0x19F6
		"--------",	-- 0x19F7
		"--------",	-- 0x19F8
		"--------",	-- 0x19F9
		"--------",	-- 0x19FA
		"--------",	-- 0x19FB
		"--------",	-- 0x19FC
		"--------",	-- 0x19FD
		"--------",	-- 0x19FE
		"--------",	-- 0x19FF
		"--------",	-- 0x1A00
		"--------",	-- 0x1A01
		"--------",	-- 0x1A02
		"--------",	-- 0x1A03
		"--------",	-- 0x1A04
		"--------",	-- 0x1A05
		"--------",	-- 0x1A06
		"--------",	-- 0x1A07
		"--------",	-- 0x1A08
		"--------",	-- 0x1A09
		"--------",	-- 0x1A0A
		"--------",	-- 0x1A0B
		"--------",	-- 0x1A0C
		"--------",	-- 0x1A0D
		"--------",	-- 0x1A0E
		"--------",	-- 0x1A0F
		"--------",	-- 0x1A10
		"--------",	-- 0x1A11
		"--------",	-- 0x1A12
		"--------",	-- 0x1A13
		"--------",	-- 0x1A14
		"--------",	-- 0x1A15
		"--------",	-- 0x1A16
		"--------",	-- 0x1A17
		"--------",	-- 0x1A18
		"--------",	-- 0x1A19
		"--------",	-- 0x1A1A
		"--------",	-- 0x1A1B
		"--------",	-- 0x1A1C
		"--------",	-- 0x1A1D
		"--------",	-- 0x1A1E
		"--------",	-- 0x1A1F
		"--------",	-- 0x1A20
		"--------",	-- 0x1A21
		"--------",	-- 0x1A22
		"--------",	-- 0x1A23
		"--------",	-- 0x1A24
		"--------",	-- 0x1A25
		"--------",	-- 0x1A26
		"--------",	-- 0x1A27
		"--------",	-- 0x1A28
		"--------",	-- 0x1A29
		"--------",	-- 0x1A2A
		"--------",	-- 0x1A2B
		"--------",	-- 0x1A2C
		"--------",	-- 0x1A2D
		"--------",	-- 0x1A2E
		"--------",	-- 0x1A2F
		"--------",	-- 0x1A30
		"--------",	-- 0x1A31
		"--------",	-- 0x1A32
		"--------",	-- 0x1A33
		"--------",	-- 0x1A34
		"--------",	-- 0x1A35
		"--------",	-- 0x1A36
		"--------",	-- 0x1A37
		"--------",	-- 0x1A38
		"--------",	-- 0x1A39
		"--------",	-- 0x1A3A
		"--------",	-- 0x1A3B
		"--------",	-- 0x1A3C
		"--------",	-- 0x1A3D
		"--------",	-- 0x1A3E
		"--------",	-- 0x1A3F
		"--------",	-- 0x1A40
		"--------",	-- 0x1A41
		"--------",	-- 0x1A42
		"--------",	-- 0x1A43
		"--------",	-- 0x1A44
		"--------",	-- 0x1A45
		"--------",	-- 0x1A46
		"--------",	-- 0x1A47
		"--------",	-- 0x1A48
		"--------",	-- 0x1A49
		"--------",	-- 0x1A4A
		"--------",	-- 0x1A4B
		"--------",	-- 0x1A4C
		"--------",	-- 0x1A4D
		"--------",	-- 0x1A4E
		"--------",	-- 0x1A4F
		"--------",	-- 0x1A50
		"--------",	-- 0x1A51
		"--------",	-- 0x1A52
		"--------",	-- 0x1A53
		"--------",	-- 0x1A54
		"--------",	-- 0x1A55
		"--------",	-- 0x1A56
		"--------",	-- 0x1A57
		"--------",	-- 0x1A58
		"--------",	-- 0x1A59
		"--------",	-- 0x1A5A
		"--------",	-- 0x1A5B
		"--------",	-- 0x1A5C
		"--------",	-- 0x1A5D
		"--------",	-- 0x1A5E
		"--------",	-- 0x1A5F
		"--------",	-- 0x1A60
		"--------",	-- 0x1A61
		"--------",	-- 0x1A62
		"--------",	-- 0x1A63
		"--------",	-- 0x1A64
		"--------",	-- 0x1A65
		"--------",	-- 0x1A66
		"--------",	-- 0x1A67
		"--------",	-- 0x1A68
		"--------",	-- 0x1A69
		"--------",	-- 0x1A6A
		"--------",	-- 0x1A6B
		"--------",	-- 0x1A6C
		"--------",	-- 0x1A6D
		"--------",	-- 0x1A6E
		"--------",	-- 0x1A6F
		"--------",	-- 0x1A70
		"--------",	-- 0x1A71
		"--------",	-- 0x1A72
		"--------",	-- 0x1A73
		"--------",	-- 0x1A74
		"--------",	-- 0x1A75
		"--------",	-- 0x1A76
		"--------",	-- 0x1A77
		"--------",	-- 0x1A78
		"--------",	-- 0x1A79
		"--------",	-- 0x1A7A
		"--------",	-- 0x1A7B
		"--------",	-- 0x1A7C
		"--------",	-- 0x1A7D
		"--------",	-- 0x1A7E
		"--------",	-- 0x1A7F
		"--------",	-- 0x1A80
		"--------",	-- 0x1A81
		"--------",	-- 0x1A82
		"--------",	-- 0x1A83
		"--------",	-- 0x1A84
		"--------",	-- 0x1A85
		"--------",	-- 0x1A86
		"--------",	-- 0x1A87
		"--------",	-- 0x1A88
		"--------",	-- 0x1A89
		"--------",	-- 0x1A8A
		"--------",	-- 0x1A8B
		"--------",	-- 0x1A8C
		"--------",	-- 0x1A8D
		"--------",	-- 0x1A8E
		"--------",	-- 0x1A8F
		"--------",	-- 0x1A90
		"--------",	-- 0x1A91
		"--------",	-- 0x1A92
		"--------",	-- 0x1A93
		"--------",	-- 0x1A94
		"--------",	-- 0x1A95
		"--------",	-- 0x1A96
		"--------",	-- 0x1A97
		"--------",	-- 0x1A98
		"--------",	-- 0x1A99
		"--------",	-- 0x1A9A
		"--------",	-- 0x1A9B
		"--------",	-- 0x1A9C
		"--------",	-- 0x1A9D
		"--------",	-- 0x1A9E
		"--------",	-- 0x1A9F
		"--------",	-- 0x1AA0
		"--------",	-- 0x1AA1
		"--------",	-- 0x1AA2
		"--------",	-- 0x1AA3
		"--------",	-- 0x1AA4
		"--------",	-- 0x1AA5
		"--------",	-- 0x1AA6
		"--------",	-- 0x1AA7
		"--------",	-- 0x1AA8
		"--------",	-- 0x1AA9
		"--------",	-- 0x1AAA
		"--------",	-- 0x1AAB
		"--------",	-- 0x1AAC
		"--------",	-- 0x1AAD
		"--------",	-- 0x1AAE
		"--------",	-- 0x1AAF
		"--------",	-- 0x1AB0
		"--------",	-- 0x1AB1
		"--------",	-- 0x1AB2
		"--------",	-- 0x1AB3
		"--------",	-- 0x1AB4
		"--------",	-- 0x1AB5
		"--------",	-- 0x1AB6
		"--------",	-- 0x1AB7
		"--------",	-- 0x1AB8
		"--------",	-- 0x1AB9
		"--------",	-- 0x1ABA
		"--------",	-- 0x1ABB
		"--------",	-- 0x1ABC
		"--------",	-- 0x1ABD
		"--------",	-- 0x1ABE
		"--------",	-- 0x1ABF
		"--------",	-- 0x1AC0
		"--------",	-- 0x1AC1
		"--------",	-- 0x1AC2
		"--------",	-- 0x1AC3
		"--------",	-- 0x1AC4
		"--------",	-- 0x1AC5
		"--------",	-- 0x1AC6
		"--------",	-- 0x1AC7
		"--------",	-- 0x1AC8
		"--------",	-- 0x1AC9
		"--------",	-- 0x1ACA
		"--------",	-- 0x1ACB
		"--------",	-- 0x1ACC
		"--------",	-- 0x1ACD
		"--------",	-- 0x1ACE
		"--------",	-- 0x1ACF
		"--------",	-- 0x1AD0
		"--------",	-- 0x1AD1
		"--------",	-- 0x1AD2
		"--------",	-- 0x1AD3
		"--------",	-- 0x1AD4
		"--------",	-- 0x1AD5
		"--------",	-- 0x1AD6
		"--------",	-- 0x1AD7
		"--------",	-- 0x1AD8
		"--------",	-- 0x1AD9
		"--------",	-- 0x1ADA
		"--------",	-- 0x1ADB
		"--------",	-- 0x1ADC
		"--------",	-- 0x1ADD
		"--------",	-- 0x1ADE
		"--------",	-- 0x1ADF
		"--------",	-- 0x1AE0
		"--------",	-- 0x1AE1
		"--------",	-- 0x1AE2
		"--------",	-- 0x1AE3
		"--------",	-- 0x1AE4
		"--------",	-- 0x1AE5
		"--------",	-- 0x1AE6
		"--------",	-- 0x1AE7
		"--------",	-- 0x1AE8
		"--------",	-- 0x1AE9
		"--------",	-- 0x1AEA
		"--------",	-- 0x1AEB
		"--------",	-- 0x1AEC
		"--------",	-- 0x1AED
		"--------",	-- 0x1AEE
		"--------",	-- 0x1AEF
		"--------",	-- 0x1AF0
		"--------",	-- 0x1AF1
		"--------",	-- 0x1AF2
		"--------",	-- 0x1AF3
		"--------",	-- 0x1AF4
		"--------",	-- 0x1AF5
		"--------",	-- 0x1AF6
		"--------",	-- 0x1AF7
		"--------",	-- 0x1AF8
		"--------",	-- 0x1AF9
		"--------",	-- 0x1AFA
		"--------",	-- 0x1AFB
		"--------",	-- 0x1AFC
		"--------",	-- 0x1AFD
		"--------",	-- 0x1AFE
		"--------",	-- 0x1AFF
		"--------",	-- 0x1B00
		"--------",	-- 0x1B01
		"--------",	-- 0x1B02
		"--------",	-- 0x1B03
		"--------",	-- 0x1B04
		"--------",	-- 0x1B05
		"--------",	-- 0x1B06
		"--------",	-- 0x1B07
		"--------",	-- 0x1B08
		"--------",	-- 0x1B09
		"--------",	-- 0x1B0A
		"--------",	-- 0x1B0B
		"--------",	-- 0x1B0C
		"--------",	-- 0x1B0D
		"--------",	-- 0x1B0E
		"--------",	-- 0x1B0F
		"--------",	-- 0x1B10
		"--------",	-- 0x1B11
		"--------",	-- 0x1B12
		"--------",	-- 0x1B13
		"--------",	-- 0x1B14
		"--------",	-- 0x1B15
		"--------",	-- 0x1B16
		"--------",	-- 0x1B17
		"--------",	-- 0x1B18
		"--------",	-- 0x1B19
		"--------",	-- 0x1B1A
		"--------",	-- 0x1B1B
		"--------",	-- 0x1B1C
		"--------",	-- 0x1B1D
		"--------",	-- 0x1B1E
		"--------",	-- 0x1B1F
		"--------",	-- 0x1B20
		"--------",	-- 0x1B21
		"--------",	-- 0x1B22
		"--------",	-- 0x1B23
		"--------",	-- 0x1B24
		"--------",	-- 0x1B25
		"--------",	-- 0x1B26
		"--------",	-- 0x1B27
		"--------",	-- 0x1B28
		"--------",	-- 0x1B29
		"--------",	-- 0x1B2A
		"--------",	-- 0x1B2B
		"--------",	-- 0x1B2C
		"--------",	-- 0x1B2D
		"--------",	-- 0x1B2E
		"--------",	-- 0x1B2F
		"--------",	-- 0x1B30
		"--------",	-- 0x1B31
		"--------",	-- 0x1B32
		"--------",	-- 0x1B33
		"--------",	-- 0x1B34
		"--------",	-- 0x1B35
		"--------",	-- 0x1B36
		"--------",	-- 0x1B37
		"--------",	-- 0x1B38
		"--------",	-- 0x1B39
		"--------",	-- 0x1B3A
		"--------",	-- 0x1B3B
		"--------",	-- 0x1B3C
		"--------",	-- 0x1B3D
		"--------",	-- 0x1B3E
		"--------",	-- 0x1B3F
		"--------",	-- 0x1B40
		"--------",	-- 0x1B41
		"--------",	-- 0x1B42
		"--------",	-- 0x1B43
		"--------",	-- 0x1B44
		"--------",	-- 0x1B45
		"--------",	-- 0x1B46
		"--------",	-- 0x1B47
		"--------",	-- 0x1B48
		"--------",	-- 0x1B49
		"--------",	-- 0x1B4A
		"--------",	-- 0x1B4B
		"--------",	-- 0x1B4C
		"--------",	-- 0x1B4D
		"--------",	-- 0x1B4E
		"--------",	-- 0x1B4F
		"--------",	-- 0x1B50
		"--------",	-- 0x1B51
		"--------",	-- 0x1B52
		"--------",	-- 0x1B53
		"--------",	-- 0x1B54
		"--------",	-- 0x1B55
		"--------",	-- 0x1B56
		"--------",	-- 0x1B57
		"--------",	-- 0x1B58
		"--------",	-- 0x1B59
		"--------",	-- 0x1B5A
		"--------",	-- 0x1B5B
		"--------",	-- 0x1B5C
		"--------",	-- 0x1B5D
		"--------",	-- 0x1B5E
		"--------",	-- 0x1B5F
		"--------",	-- 0x1B60
		"--------",	-- 0x1B61
		"--------",	-- 0x1B62
		"--------",	-- 0x1B63
		"--------",	-- 0x1B64
		"--------",	-- 0x1B65
		"--------",	-- 0x1B66
		"--------",	-- 0x1B67
		"--------",	-- 0x1B68
		"--------",	-- 0x1B69
		"--------",	-- 0x1B6A
		"--------",	-- 0x1B6B
		"--------",	-- 0x1B6C
		"--------",	-- 0x1B6D
		"--------",	-- 0x1B6E
		"--------",	-- 0x1B6F
		"--------",	-- 0x1B70
		"--------",	-- 0x1B71
		"--------",	-- 0x1B72
		"--------",	-- 0x1B73
		"--------",	-- 0x1B74
		"--------",	-- 0x1B75
		"--------",	-- 0x1B76
		"--------",	-- 0x1B77
		"--------",	-- 0x1B78
		"--------",	-- 0x1B79
		"--------",	-- 0x1B7A
		"--------",	-- 0x1B7B
		"--------",	-- 0x1B7C
		"--------",	-- 0x1B7D
		"--------",	-- 0x1B7E
		"--------",	-- 0x1B7F
		"--------",	-- 0x1B80
		"--------",	-- 0x1B81
		"--------",	-- 0x1B82
		"--------",	-- 0x1B83
		"--------",	-- 0x1B84
		"--------",	-- 0x1B85
		"--------",	-- 0x1B86
		"--------",	-- 0x1B87
		"--------",	-- 0x1B88
		"--------",	-- 0x1B89
		"--------",	-- 0x1B8A
		"--------",	-- 0x1B8B
		"--------",	-- 0x1B8C
		"--------",	-- 0x1B8D
		"--------",	-- 0x1B8E
		"--------",	-- 0x1B8F
		"--------",	-- 0x1B90
		"--------",	-- 0x1B91
		"--------",	-- 0x1B92
		"--------",	-- 0x1B93
		"--------",	-- 0x1B94
		"--------",	-- 0x1B95
		"--------",	-- 0x1B96
		"--------",	-- 0x1B97
		"--------",	-- 0x1B98
		"--------",	-- 0x1B99
		"--------",	-- 0x1B9A
		"--------",	-- 0x1B9B
		"--------",	-- 0x1B9C
		"--------",	-- 0x1B9D
		"--------",	-- 0x1B9E
		"--------",	-- 0x1B9F
		"--------",	-- 0x1BA0
		"--------",	-- 0x1BA1
		"--------",	-- 0x1BA2
		"--------",	-- 0x1BA3
		"--------",	-- 0x1BA4
		"--------",	-- 0x1BA5
		"--------",	-- 0x1BA6
		"--------",	-- 0x1BA7
		"--------",	-- 0x1BA8
		"--------",	-- 0x1BA9
		"--------",	-- 0x1BAA
		"--------",	-- 0x1BAB
		"--------",	-- 0x1BAC
		"--------",	-- 0x1BAD
		"--------",	-- 0x1BAE
		"--------",	-- 0x1BAF
		"--------",	-- 0x1BB0
		"--------",	-- 0x1BB1
		"--------",	-- 0x1BB2
		"--------",	-- 0x1BB3
		"--------",	-- 0x1BB4
		"--------",	-- 0x1BB5
		"--------",	-- 0x1BB6
		"--------",	-- 0x1BB7
		"--------",	-- 0x1BB8
		"--------",	-- 0x1BB9
		"--------",	-- 0x1BBA
		"--------",	-- 0x1BBB
		"--------",	-- 0x1BBC
		"--------",	-- 0x1BBD
		"--------",	-- 0x1BBE
		"--------",	-- 0x1BBF
		"--------",	-- 0x1BC0
		"--------",	-- 0x1BC1
		"--------",	-- 0x1BC2
		"--------",	-- 0x1BC3
		"--------",	-- 0x1BC4
		"--------",	-- 0x1BC5
		"--------",	-- 0x1BC6
		"--------",	-- 0x1BC7
		"--------",	-- 0x1BC8
		"--------",	-- 0x1BC9
		"--------",	-- 0x1BCA
		"--------",	-- 0x1BCB
		"--------",	-- 0x1BCC
		"--------",	-- 0x1BCD
		"--------",	-- 0x1BCE
		"--------",	-- 0x1BCF
		"--------",	-- 0x1BD0
		"--------",	-- 0x1BD1
		"--------",	-- 0x1BD2
		"--------",	-- 0x1BD3
		"--------",	-- 0x1BD4
		"--------",	-- 0x1BD5
		"--------",	-- 0x1BD6
		"--------",	-- 0x1BD7
		"--------",	-- 0x1BD8
		"--------",	-- 0x1BD9
		"--------",	-- 0x1BDA
		"--------",	-- 0x1BDB
		"--------",	-- 0x1BDC
		"--------",	-- 0x1BDD
		"--------",	-- 0x1BDE
		"--------",	-- 0x1BDF
		"--------",	-- 0x1BE0
		"--------",	-- 0x1BE1
		"--------",	-- 0x1BE2
		"--------",	-- 0x1BE3
		"--------",	-- 0x1BE4
		"--------",	-- 0x1BE5
		"--------",	-- 0x1BE6
		"--------",	-- 0x1BE7
		"--------",	-- 0x1BE8
		"--------",	-- 0x1BE9
		"--------",	-- 0x1BEA
		"--------",	-- 0x1BEB
		"--------",	-- 0x1BEC
		"--------",	-- 0x1BED
		"--------",	-- 0x1BEE
		"--------",	-- 0x1BEF
		"--------",	-- 0x1BF0
		"--------",	-- 0x1BF1
		"--------",	-- 0x1BF2
		"--------",	-- 0x1BF3
		"--------",	-- 0x1BF4
		"--------",	-- 0x1BF5
		"--------",	-- 0x1BF6
		"--------",	-- 0x1BF7
		"--------",	-- 0x1BF8
		"--------",	-- 0x1BF9
		"--------",	-- 0x1BFA
		"--------",	-- 0x1BFB
		"--------",	-- 0x1BFC
		"--------",	-- 0x1BFD
		"--------",	-- 0x1BFE
		"--------",	-- 0x1BFF
		"--------",	-- 0x1C00
		"--------",	-- 0x1C01
		"--------",	-- 0x1C02
		"--------",	-- 0x1C03
		"--------",	-- 0x1C04
		"--------",	-- 0x1C05
		"--------",	-- 0x1C06
		"--------",	-- 0x1C07
		"--------",	-- 0x1C08
		"--------",	-- 0x1C09
		"--------",	-- 0x1C0A
		"--------",	-- 0x1C0B
		"--------",	-- 0x1C0C
		"--------",	-- 0x1C0D
		"--------",	-- 0x1C0E
		"--------",	-- 0x1C0F
		"--------",	-- 0x1C10
		"--------",	-- 0x1C11
		"--------",	-- 0x1C12
		"--------",	-- 0x1C13
		"--------",	-- 0x1C14
		"--------",	-- 0x1C15
		"--------",	-- 0x1C16
		"--------",	-- 0x1C17
		"--------",	-- 0x1C18
		"--------",	-- 0x1C19
		"--------",	-- 0x1C1A
		"--------",	-- 0x1C1B
		"--------",	-- 0x1C1C
		"--------",	-- 0x1C1D
		"--------",	-- 0x1C1E
		"--------",	-- 0x1C1F
		"--------",	-- 0x1C20
		"--------",	-- 0x1C21
		"--------",	-- 0x1C22
		"--------",	-- 0x1C23
		"--------",	-- 0x1C24
		"--------",	-- 0x1C25
		"--------",	-- 0x1C26
		"--------",	-- 0x1C27
		"--------",	-- 0x1C28
		"--------",	-- 0x1C29
		"--------",	-- 0x1C2A
		"--------",	-- 0x1C2B
		"--------",	-- 0x1C2C
		"--------",	-- 0x1C2D
		"--------",	-- 0x1C2E
		"--------",	-- 0x1C2F
		"--------",	-- 0x1C30
		"--------",	-- 0x1C31
		"--------",	-- 0x1C32
		"--------",	-- 0x1C33
		"--------",	-- 0x1C34
		"--------",	-- 0x1C35
		"--------",	-- 0x1C36
		"--------",	-- 0x1C37
		"--------",	-- 0x1C38
		"--------",	-- 0x1C39
		"--------",	-- 0x1C3A
		"--------",	-- 0x1C3B
		"--------",	-- 0x1C3C
		"--------",	-- 0x1C3D
		"--------",	-- 0x1C3E
		"--------",	-- 0x1C3F
		"--------",	-- 0x1C40
		"--------",	-- 0x1C41
		"--------",	-- 0x1C42
		"--------",	-- 0x1C43
		"--------",	-- 0x1C44
		"--------",	-- 0x1C45
		"--------",	-- 0x1C46
		"--------",	-- 0x1C47
		"--------",	-- 0x1C48
		"--------",	-- 0x1C49
		"--------",	-- 0x1C4A
		"--------",	-- 0x1C4B
		"--------",	-- 0x1C4C
		"--------",	-- 0x1C4D
		"--------",	-- 0x1C4E
		"--------",	-- 0x1C4F
		"--------",	-- 0x1C50
		"--------",	-- 0x1C51
		"--------",	-- 0x1C52
		"--------",	-- 0x1C53
		"--------",	-- 0x1C54
		"--------",	-- 0x1C55
		"--------",	-- 0x1C56
		"--------",	-- 0x1C57
		"--------",	-- 0x1C58
		"--------",	-- 0x1C59
		"--------",	-- 0x1C5A
		"--------",	-- 0x1C5B
		"--------",	-- 0x1C5C
		"--------",	-- 0x1C5D
		"--------",	-- 0x1C5E
		"--------",	-- 0x1C5F
		"--------",	-- 0x1C60
		"--------",	-- 0x1C61
		"--------",	-- 0x1C62
		"--------",	-- 0x1C63
		"--------",	-- 0x1C64
		"--------",	-- 0x1C65
		"--------",	-- 0x1C66
		"--------",	-- 0x1C67
		"--------",	-- 0x1C68
		"--------",	-- 0x1C69
		"--------",	-- 0x1C6A
		"--------",	-- 0x1C6B
		"--------",	-- 0x1C6C
		"--------",	-- 0x1C6D
		"--------",	-- 0x1C6E
		"--------",	-- 0x1C6F
		"--------",	-- 0x1C70
		"--------",	-- 0x1C71
		"--------",	-- 0x1C72
		"--------",	-- 0x1C73
		"--------",	-- 0x1C74
		"--------",	-- 0x1C75
		"--------",	-- 0x1C76
		"--------",	-- 0x1C77
		"--------",	-- 0x1C78
		"--------",	-- 0x1C79
		"--------",	-- 0x1C7A
		"--------",	-- 0x1C7B
		"--------",	-- 0x1C7C
		"--------",	-- 0x1C7D
		"--------",	-- 0x1C7E
		"--------",	-- 0x1C7F
		"--------",	-- 0x1C80
		"--------",	-- 0x1C81
		"--------",	-- 0x1C82
		"--------",	-- 0x1C83
		"--------",	-- 0x1C84
		"--------",	-- 0x1C85
		"--------",	-- 0x1C86
		"--------",	-- 0x1C87
		"--------",	-- 0x1C88
		"--------",	-- 0x1C89
		"--------",	-- 0x1C8A
		"--------",	-- 0x1C8B
		"--------",	-- 0x1C8C
		"--------",	-- 0x1C8D
		"--------",	-- 0x1C8E
		"--------",	-- 0x1C8F
		"--------",	-- 0x1C90
		"--------",	-- 0x1C91
		"--------",	-- 0x1C92
		"--------",	-- 0x1C93
		"--------",	-- 0x1C94
		"--------",	-- 0x1C95
		"--------",	-- 0x1C96
		"--------",	-- 0x1C97
		"--------",	-- 0x1C98
		"--------",	-- 0x1C99
		"--------",	-- 0x1C9A
		"--------",	-- 0x1C9B
		"--------",	-- 0x1C9C
		"--------",	-- 0x1C9D
		"--------",	-- 0x1C9E
		"--------",	-- 0x1C9F
		"--------",	-- 0x1CA0
		"--------",	-- 0x1CA1
		"--------",	-- 0x1CA2
		"--------",	-- 0x1CA3
		"--------",	-- 0x1CA4
		"--------",	-- 0x1CA5
		"--------",	-- 0x1CA6
		"--------",	-- 0x1CA7
		"--------",	-- 0x1CA8
		"--------",	-- 0x1CA9
		"--------",	-- 0x1CAA
		"--------",	-- 0x1CAB
		"--------",	-- 0x1CAC
		"--------",	-- 0x1CAD
		"--------",	-- 0x1CAE
		"--------",	-- 0x1CAF
		"--------",	-- 0x1CB0
		"--------",	-- 0x1CB1
		"--------",	-- 0x1CB2
		"--------",	-- 0x1CB3
		"--------",	-- 0x1CB4
		"--------",	-- 0x1CB5
		"--------",	-- 0x1CB6
		"--------",	-- 0x1CB7
		"--------",	-- 0x1CB8
		"--------",	-- 0x1CB9
		"--------",	-- 0x1CBA
		"--------",	-- 0x1CBB
		"--------",	-- 0x1CBC
		"--------",	-- 0x1CBD
		"--------",	-- 0x1CBE
		"--------",	-- 0x1CBF
		"--------",	-- 0x1CC0
		"--------",	-- 0x1CC1
		"--------",	-- 0x1CC2
		"--------",	-- 0x1CC3
		"--------",	-- 0x1CC4
		"--------",	-- 0x1CC5
		"--------",	-- 0x1CC6
		"--------",	-- 0x1CC7
		"--------",	-- 0x1CC8
		"--------",	-- 0x1CC9
		"--------",	-- 0x1CCA
		"--------",	-- 0x1CCB
		"--------",	-- 0x1CCC
		"--------",	-- 0x1CCD
		"--------",	-- 0x1CCE
		"--------",	-- 0x1CCF
		"--------",	-- 0x1CD0
		"--------",	-- 0x1CD1
		"--------",	-- 0x1CD2
		"--------",	-- 0x1CD3
		"--------",	-- 0x1CD4
		"--------",	-- 0x1CD5
		"--------",	-- 0x1CD6
		"--------",	-- 0x1CD7
		"--------",	-- 0x1CD8
		"--------",	-- 0x1CD9
		"--------",	-- 0x1CDA
		"--------",	-- 0x1CDB
		"--------",	-- 0x1CDC
		"--------",	-- 0x1CDD
		"--------",	-- 0x1CDE
		"--------",	-- 0x1CDF
		"--------",	-- 0x1CE0
		"--------",	-- 0x1CE1
		"--------",	-- 0x1CE2
		"--------",	-- 0x1CE3
		"--------",	-- 0x1CE4
		"--------",	-- 0x1CE5
		"--------",	-- 0x1CE6
		"--------",	-- 0x1CE7
		"--------",	-- 0x1CE8
		"--------",	-- 0x1CE9
		"--------",	-- 0x1CEA
		"--------",	-- 0x1CEB
		"--------",	-- 0x1CEC
		"--------",	-- 0x1CED
		"--------",	-- 0x1CEE
		"--------",	-- 0x1CEF
		"--------",	-- 0x1CF0
		"--------",	-- 0x1CF1
		"--------",	-- 0x1CF2
		"--------",	-- 0x1CF3
		"--------",	-- 0x1CF4
		"--------",	-- 0x1CF5
		"--------",	-- 0x1CF6
		"--------",	-- 0x1CF7
		"--------",	-- 0x1CF8
		"--------",	-- 0x1CF9
		"--------",	-- 0x1CFA
		"--------",	-- 0x1CFB
		"--------",	-- 0x1CFC
		"--------",	-- 0x1CFD
		"--------",	-- 0x1CFE
		"--------",	-- 0x1CFF
		"--------",	-- 0x1D00
		"--------",	-- 0x1D01
		"--------",	-- 0x1D02
		"--------",	-- 0x1D03
		"--------",	-- 0x1D04
		"--------",	-- 0x1D05
		"--------",	-- 0x1D06
		"--------",	-- 0x1D07
		"--------",	-- 0x1D08
		"--------",	-- 0x1D09
		"--------",	-- 0x1D0A
		"--------",	-- 0x1D0B
		"--------",	-- 0x1D0C
		"--------",	-- 0x1D0D
		"--------",	-- 0x1D0E
		"--------",	-- 0x1D0F
		"--------",	-- 0x1D10
		"--------",	-- 0x1D11
		"--------",	-- 0x1D12
		"--------",	-- 0x1D13
		"--------",	-- 0x1D14
		"--------",	-- 0x1D15
		"--------",	-- 0x1D16
		"--------",	-- 0x1D17
		"--------",	-- 0x1D18
		"--------",	-- 0x1D19
		"--------",	-- 0x1D1A
		"--------",	-- 0x1D1B
		"--------",	-- 0x1D1C
		"--------",	-- 0x1D1D
		"--------",	-- 0x1D1E
		"--------",	-- 0x1D1F
		"--------",	-- 0x1D20
		"--------",	-- 0x1D21
		"--------",	-- 0x1D22
		"--------",	-- 0x1D23
		"--------",	-- 0x1D24
		"--------",	-- 0x1D25
		"--------",	-- 0x1D26
		"--------",	-- 0x1D27
		"--------",	-- 0x1D28
		"--------",	-- 0x1D29
		"--------",	-- 0x1D2A
		"--------",	-- 0x1D2B
		"--------",	-- 0x1D2C
		"--------",	-- 0x1D2D
		"--------",	-- 0x1D2E
		"--------",	-- 0x1D2F
		"--------",	-- 0x1D30
		"--------",	-- 0x1D31
		"--------",	-- 0x1D32
		"--------",	-- 0x1D33
		"--------",	-- 0x1D34
		"--------",	-- 0x1D35
		"--------",	-- 0x1D36
		"--------",	-- 0x1D37
		"--------",	-- 0x1D38
		"--------",	-- 0x1D39
		"--------",	-- 0x1D3A
		"--------",	-- 0x1D3B
		"--------",	-- 0x1D3C
		"--------",	-- 0x1D3D
		"--------",	-- 0x1D3E
		"--------",	-- 0x1D3F
		"--------",	-- 0x1D40
		"--------",	-- 0x1D41
		"--------",	-- 0x1D42
		"--------",	-- 0x1D43
		"--------",	-- 0x1D44
		"--------",	-- 0x1D45
		"--------",	-- 0x1D46
		"--------",	-- 0x1D47
		"--------",	-- 0x1D48
		"--------",	-- 0x1D49
		"--------",	-- 0x1D4A
		"--------",	-- 0x1D4B
		"--------",	-- 0x1D4C
		"--------",	-- 0x1D4D
		"--------",	-- 0x1D4E
		"--------",	-- 0x1D4F
		"--------",	-- 0x1D50
		"--------",	-- 0x1D51
		"--------",	-- 0x1D52
		"--------",	-- 0x1D53
		"--------",	-- 0x1D54
		"--------",	-- 0x1D55
		"--------",	-- 0x1D56
		"--------",	-- 0x1D57
		"--------",	-- 0x1D58
		"--------",	-- 0x1D59
		"--------",	-- 0x1D5A
		"--------",	-- 0x1D5B
		"--------",	-- 0x1D5C
		"--------",	-- 0x1D5D
		"--------",	-- 0x1D5E
		"--------",	-- 0x1D5F
		"--------",	-- 0x1D60
		"--------",	-- 0x1D61
		"--------",	-- 0x1D62
		"--------",	-- 0x1D63
		"--------",	-- 0x1D64
		"--------",	-- 0x1D65
		"--------",	-- 0x1D66
		"--------",	-- 0x1D67
		"--------",	-- 0x1D68
		"--------",	-- 0x1D69
		"--------",	-- 0x1D6A
		"--------",	-- 0x1D6B
		"--------",	-- 0x1D6C
		"--------",	-- 0x1D6D
		"--------",	-- 0x1D6E
		"--------",	-- 0x1D6F
		"--------",	-- 0x1D70
		"--------",	-- 0x1D71
		"--------",	-- 0x1D72
		"--------",	-- 0x1D73
		"--------",	-- 0x1D74
		"--------",	-- 0x1D75
		"--------",	-- 0x1D76
		"--------",	-- 0x1D77
		"--------",	-- 0x1D78
		"--------",	-- 0x1D79
		"--------",	-- 0x1D7A
		"--------",	-- 0x1D7B
		"--------",	-- 0x1D7C
		"--------",	-- 0x1D7D
		"--------",	-- 0x1D7E
		"--------",	-- 0x1D7F
		"--------",	-- 0x1D80
		"--------",	-- 0x1D81
		"--------",	-- 0x1D82
		"--------",	-- 0x1D83
		"--------",	-- 0x1D84
		"--------",	-- 0x1D85
		"--------",	-- 0x1D86
		"--------",	-- 0x1D87
		"--------",	-- 0x1D88
		"--------",	-- 0x1D89
		"--------",	-- 0x1D8A
		"--------",	-- 0x1D8B
		"--------",	-- 0x1D8C
		"--------",	-- 0x1D8D
		"--------",	-- 0x1D8E
		"--------",	-- 0x1D8F
		"--------",	-- 0x1D90
		"--------",	-- 0x1D91
		"--------",	-- 0x1D92
		"--------",	-- 0x1D93
		"--------",	-- 0x1D94
		"--------",	-- 0x1D95
		"--------",	-- 0x1D96
		"--------",	-- 0x1D97
		"--------",	-- 0x1D98
		"--------",	-- 0x1D99
		"--------",	-- 0x1D9A
		"--------",	-- 0x1D9B
		"--------",	-- 0x1D9C
		"--------",	-- 0x1D9D
		"--------",	-- 0x1D9E
		"--------",	-- 0x1D9F
		"--------",	-- 0x1DA0
		"--------",	-- 0x1DA1
		"--------",	-- 0x1DA2
		"--------",	-- 0x1DA3
		"--------",	-- 0x1DA4
		"--------",	-- 0x1DA5
		"--------",	-- 0x1DA6
		"--------",	-- 0x1DA7
		"--------",	-- 0x1DA8
		"--------",	-- 0x1DA9
		"--------",	-- 0x1DAA
		"--------",	-- 0x1DAB
		"--------",	-- 0x1DAC
		"--------",	-- 0x1DAD
		"--------",	-- 0x1DAE
		"--------",	-- 0x1DAF
		"--------",	-- 0x1DB0
		"--------",	-- 0x1DB1
		"--------",	-- 0x1DB2
		"--------",	-- 0x1DB3
		"--------",	-- 0x1DB4
		"--------",	-- 0x1DB5
		"--------",	-- 0x1DB6
		"--------",	-- 0x1DB7
		"--------",	-- 0x1DB8
		"--------",	-- 0x1DB9
		"--------",	-- 0x1DBA
		"--------",	-- 0x1DBB
		"--------",	-- 0x1DBC
		"--------",	-- 0x1DBD
		"--------",	-- 0x1DBE
		"--------",	-- 0x1DBF
		"--------",	-- 0x1DC0
		"--------",	-- 0x1DC1
		"--------",	-- 0x1DC2
		"--------",	-- 0x1DC3
		"--------",	-- 0x1DC4
		"--------",	-- 0x1DC5
		"--------",	-- 0x1DC6
		"--------",	-- 0x1DC7
		"--------",	-- 0x1DC8
		"--------",	-- 0x1DC9
		"--------",	-- 0x1DCA
		"--------",	-- 0x1DCB
		"--------",	-- 0x1DCC
		"--------",	-- 0x1DCD
		"--------",	-- 0x1DCE
		"--------",	-- 0x1DCF
		"--------",	-- 0x1DD0
		"--------",	-- 0x1DD1
		"--------",	-- 0x1DD2
		"--------",	-- 0x1DD3
		"--------",	-- 0x1DD4
		"--------",	-- 0x1DD5
		"--------",	-- 0x1DD6
		"--------",	-- 0x1DD7
		"--------",	-- 0x1DD8
		"--------",	-- 0x1DD9
		"--------",	-- 0x1DDA
		"--------",	-- 0x1DDB
		"--------",	-- 0x1DDC
		"--------",	-- 0x1DDD
		"--------",	-- 0x1DDE
		"--------",	-- 0x1DDF
		"--------",	-- 0x1DE0
		"--------",	-- 0x1DE1
		"--------",	-- 0x1DE2
		"--------",	-- 0x1DE3
		"--------",	-- 0x1DE4
		"--------",	-- 0x1DE5
		"--------",	-- 0x1DE6
		"--------",	-- 0x1DE7
		"--------",	-- 0x1DE8
		"--------",	-- 0x1DE9
		"--------",	-- 0x1DEA
		"--------",	-- 0x1DEB
		"--------",	-- 0x1DEC
		"--------",	-- 0x1DED
		"--------",	-- 0x1DEE
		"--------",	-- 0x1DEF
		"--------",	-- 0x1DF0
		"--------",	-- 0x1DF1
		"--------",	-- 0x1DF2
		"--------",	-- 0x1DF3
		"--------",	-- 0x1DF4
		"--------",	-- 0x1DF5
		"--------",	-- 0x1DF6
		"--------",	-- 0x1DF7
		"--------",	-- 0x1DF8
		"--------",	-- 0x1DF9
		"--------",	-- 0x1DFA
		"--------",	-- 0x1DFB
		"--------",	-- 0x1DFC
		"--------",	-- 0x1DFD
		"--------",	-- 0x1DFE
		"--------",	-- 0x1DFF
		"--------",	-- 0x1E00
		"--------",	-- 0x1E01
		"--------",	-- 0x1E02
		"--------",	-- 0x1E03
		"--------",	-- 0x1E04
		"--------",	-- 0x1E05
		"--------",	-- 0x1E06
		"--------",	-- 0x1E07
		"--------",	-- 0x1E08
		"--------",	-- 0x1E09
		"--------",	-- 0x1E0A
		"--------",	-- 0x1E0B
		"--------",	-- 0x1E0C
		"--------",	-- 0x1E0D
		"--------",	-- 0x1E0E
		"--------",	-- 0x1E0F
		"--------",	-- 0x1E10
		"--------",	-- 0x1E11
		"--------",	-- 0x1E12
		"--------",	-- 0x1E13
		"--------",	-- 0x1E14
		"--------",	-- 0x1E15
		"--------",	-- 0x1E16
		"--------",	-- 0x1E17
		"--------",	-- 0x1E18
		"--------",	-- 0x1E19
		"--------",	-- 0x1E1A
		"--------",	-- 0x1E1B
		"--------",	-- 0x1E1C
		"--------",	-- 0x1E1D
		"--------",	-- 0x1E1E
		"--------",	-- 0x1E1F
		"--------",	-- 0x1E20
		"--------",	-- 0x1E21
		"--------",	-- 0x1E22
		"--------",	-- 0x1E23
		"--------",	-- 0x1E24
		"--------",	-- 0x1E25
		"--------",	-- 0x1E26
		"--------",	-- 0x1E27
		"--------",	-- 0x1E28
		"--------",	-- 0x1E29
		"--------",	-- 0x1E2A
		"--------",	-- 0x1E2B
		"--------",	-- 0x1E2C
		"--------",	-- 0x1E2D
		"--------",	-- 0x1E2E
		"--------",	-- 0x1E2F
		"--------",	-- 0x1E30
		"--------",	-- 0x1E31
		"--------",	-- 0x1E32
		"--------",	-- 0x1E33
		"--------",	-- 0x1E34
		"--------",	-- 0x1E35
		"--------",	-- 0x1E36
		"--------",	-- 0x1E37
		"--------",	-- 0x1E38
		"--------",	-- 0x1E39
		"--------",	-- 0x1E3A
		"--------",	-- 0x1E3B
		"--------",	-- 0x1E3C
		"--------",	-- 0x1E3D
		"--------",	-- 0x1E3E
		"--------",	-- 0x1E3F
		"--------",	-- 0x1E40
		"--------",	-- 0x1E41
		"--------",	-- 0x1E42
		"--------",	-- 0x1E43
		"--------",	-- 0x1E44
		"--------",	-- 0x1E45
		"--------",	-- 0x1E46
		"--------",	-- 0x1E47
		"--------",	-- 0x1E48
		"--------",	-- 0x1E49
		"--------",	-- 0x1E4A
		"--------",	-- 0x1E4B
		"--------",	-- 0x1E4C
		"--------",	-- 0x1E4D
		"--------",	-- 0x1E4E
		"--------",	-- 0x1E4F
		"--------",	-- 0x1E50
		"--------",	-- 0x1E51
		"--------",	-- 0x1E52
		"--------",	-- 0x1E53
		"--------",	-- 0x1E54
		"--------",	-- 0x1E55
		"--------",	-- 0x1E56
		"--------",	-- 0x1E57
		"--------",	-- 0x1E58
		"--------",	-- 0x1E59
		"--------",	-- 0x1E5A
		"--------",	-- 0x1E5B
		"--------",	-- 0x1E5C
		"--------",	-- 0x1E5D
		"--------",	-- 0x1E5E
		"--------",	-- 0x1E5F
		"--------",	-- 0x1E60
		"--------",	-- 0x1E61
		"--------",	-- 0x1E62
		"--------",	-- 0x1E63
		"--------",	-- 0x1E64
		"--------",	-- 0x1E65
		"--------",	-- 0x1E66
		"--------",	-- 0x1E67
		"--------",	-- 0x1E68
		"--------",	-- 0x1E69
		"--------",	-- 0x1E6A
		"--------",	-- 0x1E6B
		"--------",	-- 0x1E6C
		"--------",	-- 0x1E6D
		"--------",	-- 0x1E6E
		"--------",	-- 0x1E6F
		"--------",	-- 0x1E70
		"--------",	-- 0x1E71
		"--------",	-- 0x1E72
		"--------",	-- 0x1E73
		"--------",	-- 0x1E74
		"--------",	-- 0x1E75
		"--------",	-- 0x1E76
		"--------",	-- 0x1E77
		"--------",	-- 0x1E78
		"--------",	-- 0x1E79
		"--------",	-- 0x1E7A
		"--------",	-- 0x1E7B
		"--------",	-- 0x1E7C
		"--------",	-- 0x1E7D
		"--------",	-- 0x1E7E
		"--------",	-- 0x1E7F
		"--------",	-- 0x1E80
		"--------",	-- 0x1E81
		"--------",	-- 0x1E82
		"--------",	-- 0x1E83
		"--------",	-- 0x1E84
		"--------",	-- 0x1E85
		"--------",	-- 0x1E86
		"--------",	-- 0x1E87
		"--------",	-- 0x1E88
		"--------",	-- 0x1E89
		"--------",	-- 0x1E8A
		"--------",	-- 0x1E8B
		"--------",	-- 0x1E8C
		"--------",	-- 0x1E8D
		"--------",	-- 0x1E8E
		"--------",	-- 0x1E8F
		"--------",	-- 0x1E90
		"--------",	-- 0x1E91
		"--------",	-- 0x1E92
		"--------",	-- 0x1E93
		"--------",	-- 0x1E94
		"--------",	-- 0x1E95
		"--------",	-- 0x1E96
		"--------",	-- 0x1E97
		"--------",	-- 0x1E98
		"--------",	-- 0x1E99
		"--------",	-- 0x1E9A
		"--------",	-- 0x1E9B
		"--------",	-- 0x1E9C
		"--------",	-- 0x1E9D
		"--------",	-- 0x1E9E
		"--------",	-- 0x1E9F
		"--------",	-- 0x1EA0
		"--------",	-- 0x1EA1
		"--------",	-- 0x1EA2
		"--------",	-- 0x1EA3
		"--------",	-- 0x1EA4
		"--------",	-- 0x1EA5
		"--------",	-- 0x1EA6
		"--------",	-- 0x1EA7
		"--------",	-- 0x1EA8
		"--------",	-- 0x1EA9
		"--------",	-- 0x1EAA
		"--------",	-- 0x1EAB
		"--------",	-- 0x1EAC
		"--------",	-- 0x1EAD
		"--------",	-- 0x1EAE
		"--------",	-- 0x1EAF
		"--------",	-- 0x1EB0
		"--------",	-- 0x1EB1
		"--------",	-- 0x1EB2
		"--------",	-- 0x1EB3
		"--------",	-- 0x1EB4
		"--------",	-- 0x1EB5
		"--------",	-- 0x1EB6
		"--------",	-- 0x1EB7
		"--------",	-- 0x1EB8
		"--------",	-- 0x1EB9
		"--------",	-- 0x1EBA
		"--------",	-- 0x1EBB
		"--------",	-- 0x1EBC
		"--------",	-- 0x1EBD
		"--------",	-- 0x1EBE
		"--------",	-- 0x1EBF
		"--------",	-- 0x1EC0
		"--------",	-- 0x1EC1
		"--------",	-- 0x1EC2
		"--------",	-- 0x1EC3
		"--------",	-- 0x1EC4
		"--------",	-- 0x1EC5
		"--------",	-- 0x1EC6
		"--------",	-- 0x1EC7
		"--------",	-- 0x1EC8
		"--------",	-- 0x1EC9
		"--------",	-- 0x1ECA
		"--------",	-- 0x1ECB
		"--------",	-- 0x1ECC
		"--------",	-- 0x1ECD
		"--------",	-- 0x1ECE
		"--------",	-- 0x1ECF
		"--------",	-- 0x1ED0
		"--------",	-- 0x1ED1
		"--------",	-- 0x1ED2
		"--------",	-- 0x1ED3
		"--------",	-- 0x1ED4
		"--------",	-- 0x1ED5
		"--------",	-- 0x1ED6
		"--------",	-- 0x1ED7
		"--------",	-- 0x1ED8
		"--------",	-- 0x1ED9
		"--------",	-- 0x1EDA
		"--------",	-- 0x1EDB
		"--------",	-- 0x1EDC
		"--------",	-- 0x1EDD
		"--------",	-- 0x1EDE
		"--------",	-- 0x1EDF
		"--------",	-- 0x1EE0
		"--------",	-- 0x1EE1
		"--------",	-- 0x1EE2
		"--------",	-- 0x1EE3
		"--------",	-- 0x1EE4
		"--------",	-- 0x1EE5
		"--------",	-- 0x1EE6
		"--------",	-- 0x1EE7
		"--------",	-- 0x1EE8
		"--------",	-- 0x1EE9
		"--------",	-- 0x1EEA
		"--------",	-- 0x1EEB
		"--------",	-- 0x1EEC
		"--------",	-- 0x1EED
		"--------",	-- 0x1EEE
		"--------",	-- 0x1EEF
		"--------",	-- 0x1EF0
		"--------",	-- 0x1EF1
		"--------",	-- 0x1EF2
		"--------",	-- 0x1EF3
		"--------",	-- 0x1EF4
		"--------",	-- 0x1EF5
		"--------",	-- 0x1EF6
		"--------",	-- 0x1EF7
		"--------",	-- 0x1EF8
		"--------",	-- 0x1EF9
		"--------",	-- 0x1EFA
		"--------",	-- 0x1EFB
		"--------",	-- 0x1EFC
		"--------",	-- 0x1EFD
		"--------",	-- 0x1EFE
		"--------",	-- 0x1EFF
		"--------",	-- 0x1F00
		"--------",	-- 0x1F01
		"--------",	-- 0x1F02
		"--------",	-- 0x1F03
		"--------",	-- 0x1F04
		"--------",	-- 0x1F05
		"--------",	-- 0x1F06
		"--------",	-- 0x1F07
		"--------",	-- 0x1F08
		"--------",	-- 0x1F09
		"--------",	-- 0x1F0A
		"--------",	-- 0x1F0B
		"--------",	-- 0x1F0C
		"--------",	-- 0x1F0D
		"--------",	-- 0x1F0E
		"--------",	-- 0x1F0F
		"--------",	-- 0x1F10
		"--------",	-- 0x1F11
		"--------",	-- 0x1F12
		"--------",	-- 0x1F13
		"--------",	-- 0x1F14
		"--------",	-- 0x1F15
		"--------",	-- 0x1F16
		"--------",	-- 0x1F17
		"--------",	-- 0x1F18
		"--------",	-- 0x1F19
		"--------",	-- 0x1F1A
		"--------",	-- 0x1F1B
		"--------",	-- 0x1F1C
		"--------",	-- 0x1F1D
		"--------",	-- 0x1F1E
		"--------",	-- 0x1F1F
		"--------",	-- 0x1F20
		"--------",	-- 0x1F21
		"--------",	-- 0x1F22
		"--------",	-- 0x1F23
		"--------",	-- 0x1F24
		"--------",	-- 0x1F25
		"--------",	-- 0x1F26
		"--------",	-- 0x1F27
		"--------",	-- 0x1F28
		"--------",	-- 0x1F29
		"--------",	-- 0x1F2A
		"--------",	-- 0x1F2B
		"--------",	-- 0x1F2C
		"--------",	-- 0x1F2D
		"--------",	-- 0x1F2E
		"--------",	-- 0x1F2F
		"--------",	-- 0x1F30
		"--------",	-- 0x1F31
		"--------",	-- 0x1F32
		"--------",	-- 0x1F33
		"--------",	-- 0x1F34
		"--------",	-- 0x1F35
		"--------",	-- 0x1F36
		"--------",	-- 0x1F37
		"--------",	-- 0x1F38
		"--------",	-- 0x1F39
		"--------",	-- 0x1F3A
		"--------",	-- 0x1F3B
		"--------",	-- 0x1F3C
		"--------",	-- 0x1F3D
		"--------",	-- 0x1F3E
		"--------",	-- 0x1F3F
		"--------",	-- 0x1F40
		"--------",	-- 0x1F41
		"--------",	-- 0x1F42
		"--------",	-- 0x1F43
		"--------",	-- 0x1F44
		"--------",	-- 0x1F45
		"--------",	-- 0x1F46
		"--------",	-- 0x1F47
		"--------",	-- 0x1F48
		"--------",	-- 0x1F49
		"--------",	-- 0x1F4A
		"--------",	-- 0x1F4B
		"--------",	-- 0x1F4C
		"--------",	-- 0x1F4D
		"--------",	-- 0x1F4E
		"--------",	-- 0x1F4F
		"--------",	-- 0x1F50
		"--------",	-- 0x1F51
		"--------",	-- 0x1F52
		"--------",	-- 0x1F53
		"--------",	-- 0x1F54
		"--------",	-- 0x1F55
		"--------",	-- 0x1F56
		"--------",	-- 0x1F57
		"--------",	-- 0x1F58
		"--------",	-- 0x1F59
		"--------",	-- 0x1F5A
		"--------",	-- 0x1F5B
		"--------",	-- 0x1F5C
		"--------",	-- 0x1F5D
		"--------",	-- 0x1F5E
		"--------",	-- 0x1F5F
		"--------",	-- 0x1F60
		"--------",	-- 0x1F61
		"--------",	-- 0x1F62
		"--------",	-- 0x1F63
		"--------",	-- 0x1F64
		"--------",	-- 0x1F65
		"--------",	-- 0x1F66
		"--------",	-- 0x1F67
		"--------",	-- 0x1F68
		"--------",	-- 0x1F69
		"--------",	-- 0x1F6A
		"--------",	-- 0x1F6B
		"--------",	-- 0x1F6C
		"--------",	-- 0x1F6D
		"--------",	-- 0x1F6E
		"--------",	-- 0x1F6F
		"--------",	-- 0x1F70
		"--------",	-- 0x1F71
		"--------",	-- 0x1F72
		"--------",	-- 0x1F73
		"--------",	-- 0x1F74
		"--------",	-- 0x1F75
		"--------",	-- 0x1F76
		"--------",	-- 0x1F77
		"--------",	-- 0x1F78
		"--------",	-- 0x1F79
		"--------",	-- 0x1F7A
		"--------",	-- 0x1F7B
		"--------",	-- 0x1F7C
		"--------",	-- 0x1F7D
		"--------",	-- 0x1F7E
		"--------",	-- 0x1F7F
		"--------",	-- 0x1F80
		"--------",	-- 0x1F81
		"--------",	-- 0x1F82
		"--------",	-- 0x1F83
		"--------",	-- 0x1F84
		"--------",	-- 0x1F85
		"--------",	-- 0x1F86
		"--------",	-- 0x1F87
		"--------",	-- 0x1F88
		"--------",	-- 0x1F89
		"--------",	-- 0x1F8A
		"--------",	-- 0x1F8B
		"--------",	-- 0x1F8C
		"--------",	-- 0x1F8D
		"--------",	-- 0x1F8E
		"--------",	-- 0x1F8F
		"--------",	-- 0x1F90
		"--------",	-- 0x1F91
		"--------",	-- 0x1F92
		"--------",	-- 0x1F93
		"--------",	-- 0x1F94
		"--------",	-- 0x1F95
		"--------",	-- 0x1F96
		"--------",	-- 0x1F97
		"--------",	-- 0x1F98
		"--------",	-- 0x1F99
		"--------",	-- 0x1F9A
		"--------",	-- 0x1F9B
		"--------",	-- 0x1F9C
		"--------",	-- 0x1F9D
		"--------",	-- 0x1F9E
		"--------",	-- 0x1F9F
		"--------",	-- 0x1FA0
		"--------",	-- 0x1FA1
		"--------",	-- 0x1FA2
		"--------",	-- 0x1FA3
		"--------",	-- 0x1FA4
		"--------",	-- 0x1FA5
		"--------",	-- 0x1FA6
		"--------",	-- 0x1FA7
		"--------",	-- 0x1FA8
		"--------",	-- 0x1FA9
		"--------",	-- 0x1FAA
		"--------",	-- 0x1FAB
		"--------",	-- 0x1FAC
		"--------",	-- 0x1FAD
		"--------",	-- 0x1FAE
		"--------",	-- 0x1FAF
		"--------",	-- 0x1FB0
		"--------",	-- 0x1FB1
		"--------",	-- 0x1FB2
		"--------",	-- 0x1FB3
		"--------",	-- 0x1FB4
		"--------",	-- 0x1FB5
		"--------",	-- 0x1FB6
		"--------",	-- 0x1FB7
		"--------",	-- 0x1FB8
		"--------",	-- 0x1FB9
		"--------",	-- 0x1FBA
		"--------",	-- 0x1FBB
		"--------",	-- 0x1FBC
		"--------",	-- 0x1FBD
		"--------",	-- 0x1FBE
		"--------",	-- 0x1FBF
		"--------",	-- 0x1FC0
		"--------",	-- 0x1FC1
		"--------",	-- 0x1FC2
		"--------",	-- 0x1FC3
		"--------",	-- 0x1FC4
		"--------",	-- 0x1FC5
		"--------",	-- 0x1FC6
		"--------",	-- 0x1FC7
		"--------",	-- 0x1FC8
		"--------",	-- 0x1FC9
		"--------",	-- 0x1FCA
		"--------",	-- 0x1FCB
		"--------",	-- 0x1FCC
		"--------",	-- 0x1FCD
		"--------",	-- 0x1FCE
		"--------",	-- 0x1FCF
		"--------",	-- 0x1FD0
		"--------",	-- 0x1FD1
		"--------",	-- 0x1FD2
		"--------",	-- 0x1FD3
		"--------",	-- 0x1FD4
		"--------",	-- 0x1FD5
		"--------",	-- 0x1FD6
		"--------",	-- 0x1FD7
		"--------",	-- 0x1FD8
		"--------",	-- 0x1FD9
		"--------",	-- 0x1FDA
		"--------",	-- 0x1FDB
		"--------",	-- 0x1FDC
		"--------",	-- 0x1FDD
		"--------",	-- 0x1FDE
		"--------",	-- 0x1FDF
		"--------",	-- 0x1FE0
		"--------",	-- 0x1FE1
		"--------",	-- 0x1FE2
		"--------",	-- 0x1FE3
		"--------",	-- 0x1FE4
		"--------",	-- 0x1FE5
		"--------",	-- 0x1FE6
		"--------",	-- 0x1FE7
		"--------",	-- 0x1FE8
		"--------",	-- 0x1FE9
		"--------",	-- 0x1FEA
		"--------",	-- 0x1FEB
		"--------",	-- 0x1FEC
		"--------",	-- 0x1FED
		"--------",	-- 0x1FEE
		"--------",	-- 0x1FEF
		"--------",	-- 0x1FF0
		"--------",	-- 0x1FF1
		"--------",	-- 0x1FF2
		"--------",	-- 0x1FF3
		"--------",	-- 0x1FF4
		"--------",	-- 0x1FF5
		"--------",	-- 0x1FF6
		"--------",	-- 0x1FF7
		"--------",	-- 0x1FF8
		"--------",	-- 0x1FF9
		"--------",	-- 0x1FFA
		"--------",	-- 0x1FFB
		"--------",	-- 0x1FFC
		"--------",	-- 0x1FFD
		"--------",	-- 0x1FFE
		"--------");	-- 0x1FFF
begin
	D <= ROM(to_integer(unsigned(A))) when CE_n = '0' and OE_n = '0' else (others => 'Z');
end;
